* SPICE NETLIST
***************************************

.SUBCKT L POS NEG SUB
.ENDS
***************************************
.SUBCKT ICV_1
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT YA2GSD O E2 E8 E4 I SR E
** N=8 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_2 1 2 3 4 5
** N=6 EP=5 IP=8 FDC=0
X0 1 2 2 2 3 2 4 YA2GSD $T=1411120 1155550 0 90 $X=1271620 $Y=1158400
.ENDS
***************************************
.SUBCKT ICV_3 1 2 3 4 5 6 7 8
** N=10 EP=8 IP=16 FDC=0
X0 6 2 2 2 1 2 5 YA2GSD $T=1411120 939930 0 90 $X=1271620 $Y=942780
X1 7 3 3 3 4 3 5 YA2GSD $T=1411120 1047740 0 90 $X=1271620 $Y=1050590
.ENDS
***************************************
.SUBCKT ICV_4 1 2 3 4 7
** N=20 EP=5 IP=8 FDC=0
X0 3 1 1 1 2 1 4 YA2GSD $T=1411120 832130 0 90 $X=1271620 $Y=834980
.ENDS
***************************************
.SUBCKT ICV_5 1 2 3 4 5 6 7 8 10
** N=11 EP=9 IP=16 FDC=0
X0 6 1 1 1 7 2 3 YA2GSD $T=1411120 400930 0 90 $X=1271620 $Y=403780
X1 8 2 2 2 4 2 5 YA2GSD $T=1411120 508730 0 90 $X=1271620 $Y=511580
.ENDS
***************************************
.SUBCKT ICV_6 1 2 3 4 5 6 7 8 9
** N=11 EP=9 IP=16 FDC=0
X0 5 1 1 1 2 4 3 YA2GSD $T=1411120 185310 0 90 $X=1271620 $Y=188160
X1 6 4 4 4 7 8 3 YA2GSD $T=1411120 293120 0 90 $X=1271620 $Y=295970
.ENDS
***************************************
.SUBCKT ICV_7
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT XMD I SMT PU PD O
** N=6 EP=5 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_8 1 2 3 4 5 6 9
** N=11 EP=7 IP=12 FDC=0
X0 2 1 1 1 3 XMD $T=1150000 1403480 0 180 $X=1090230 $Y=1263980
X1 4 5 1 1 6 XMD $T=1241810 1403480 0 180 $X=1182040 $Y=1263980
.ENDS
***************************************
.SUBCKT INV1S I VCC O GND
** N=5 EP=4 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT BUF1 I VCC GND O
** N=5 EP=4 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_9 1 2 3 4 5 10
** N=10 EP=6 IP=10 FDC=0
X0 2 5 3 1 INV1S $T=1114760 1183280 1 0 $X=1114760 $Y=1177860
X1 3 5 1 4 BUF1 $T=1178000 1183280 1 0 $X=1178000 $Y=1177860
.ENDS
***************************************
.SUBCKT ICV_10 1 2 3 4 7 9
** N=9 EP=6 IP=10 FDC=0
X0 2 1 7 4 BUF1 $T=1183580 981680 1 0 $X=1183580 $Y=976260
X1 3 1 7 2 BUF1 $T=1183580 1092560 1 0 $X=1183580 $Y=1087140
.ENDS
***************************************
.SUBCKT ICV_11 1 2 3 4 7
** N=7 EP=5 IP=5 FDC=0
X0 1 3 4 2 BUF1 $T=1183580 890960 1 0 $X=1183580 $Y=885540
.ENDS
***************************************
.SUBCKT TIE1 O VCC GND
** N=4 EP=3 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_12 1 2 3 4 6 7 9
** N=10 EP=7 IP=19 FDC=0
X0 1 6 7 2 BUF1 $T=1182340 427280 1 0 $X=1182340 $Y=421860
X1 10 6 7 3 BUF1 $T=1184200 437360 0 0 $X=1184200 $Y=436980
X2 10 6 7 4 BUF1 $T=1184200 528080 0 0 $X=1184200 $Y=527700
X3 10 6 7 TIE1 $T=1184820 518000 0 0 $X=1184820 $Y=517620
.ENDS
***************************************
.SUBCKT ICV_13 2 3 4 5 6 7 8 9 10 14
** N=14 EP=10 IP=25 FDC=0
X0 3 2 10 4 BUF1 $T=1068260 225680 1 0 $X=1068260 $Y=220260
X1 6 2 10 5 BUF1 $T=1088720 225680 0 180 $X=1086240 $Y=220260
X2 4 2 10 7 BUF1 $T=1179860 225680 1 0 $X=1179860 $Y=220260
X3 7 2 10 8 BUF1 $T=1181720 235760 1 0 $X=1181720 $Y=230340
X4 8 2 10 9 BUF1 $T=1182960 316400 0 0 $X=1182960 $Y=316020
.ENDS
***************************************
.SUBCKT ICV_14 1 2 3 4 5 6 7 8 10
** N=11 EP=9 IP=16 FDC=0
X0 3 1 4 4 5 4 2 YA2GSD $T=1054000 0 0 0 $X=1056850 $Y=0
X1 6 4 4 7 8 7 2 YA2GSD $T=1162500 0 0 0 $X=1165350 $Y=0
.ENDS
***************************************
.SUBCKT ICV_15 1 2 3 4 5 6 7 8 9 10 13
** N=14 EP=11 IP=18 FDC=0
X0 3 1 1 4 5 XMD $T=874570 1403480 0 180 $X=814800 $Y=1263980
X1 6 2 2 2 7 XMD $T=966380 1403480 0 180 $X=906610 $Y=1263980
X2 8 9 2 2 10 XMD $T=1058190 1403480 0 180 $X=998420 $Y=1263980
.ENDS
***************************************
.SUBCKT ICV_16 1 2 3 4 5 6 7 14
** N=14 EP=8 IP=20 FDC=0
X0 4 7 5 1 INV1S $T=1026720 1183280 1 0 $X=1026720 $Y=1177860
X1 5 7 6 1 INV1S $T=1038500 1183280 0 180 $X=1037260 $Y=1177860
X2 3 7 1 2 BUF1 $T=841960 1183280 0 180 $X=839480 $Y=1177860
X3 3 7 1 4 BUF1 $T=930000 1183280 1 0 $X=930000 $Y=1177860
.ENDS
***************************************
.SUBCKT ICV_17
** N=6 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT TIE0 O VCC GND
** N=4 EP=3 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_18 2 3 4 5 6
** N=6 EP=5 IP=9 FDC=0
X0 3 4 2 5 INV1S $T=846300 780080 1 180 $X=845060 $Y=779700
X1 3 4 5 TIE0 $T=847540 800240 1 0 $X=847540 $Y=794820
.ENDS
***************************************
.SUBCKT ICV_19
** N=6 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_20 2 3 4 5 7 13
** N=13 EP=6 IP=10 FDC=0
X0 3 2 4 7 INV1S $T=848780 225680 1 0 $X=848780 $Y=220260
X1 4 2 7 5 BUF1 $T=903960 225680 1 0 $X=903960 $Y=220260
.ENDS
***************************************
.SUBCKT ICV_21 1 2 3 4 5 6 7 10
** N=12 EP=8 IP=16 FDC=0
X0 3 1 1 1 4 1 5 YA2GSD $T=837000 0 0 0 $X=839850 $Y=0
X1 6 2 2 2 7 2 5 YA2GSD $T=945500 0 0 0 $X=948350 $Y=0
.ENDS
***************************************
.SUBCKT ICV_22 1 2 3 10 11 12 13 14 15 39
** N=53 EP=10 IP=18 FDC=0
X0 10 2 1 1 11 XMD $T=415550 1403480 0 180 $X=355780 $Y=1263980
X1 12 2 2 2 13 XMD $T=507360 1403480 0 180 $X=447590 $Y=1263980
X2 14 3 3 2 15 XMD $T=599170 1403480 0 180 $X=539400 $Y=1263980
.ENDS
***************************************
.SUBCKT ICV_23 1 2 3 7 14 41
** N=41 EP=6 IP=10 FDC=0
X0 3 14 1 2 BUF1 $T=389360 1183280 0 180 $X=386880 $Y=1177860
X1 7 14 1 3 BUF1 $T=570400 1183280 0 180 $X=567920 $Y=1177860
.ENDS
***************************************
.SUBCKT ICV_24
** N=19 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT QDFFRBN D CK RB VCC GND Q
** N=7 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AOI22S A1 B1 O B2 GND A2 VCC
** N=8 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ND2 I1 O I2 GND VCC
** N=6 EP=5 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT FA1S CO VCC A B CI GND S
** N=8 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT NR2 I1 VCC O I2 GND
** N=6 EP=5 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT HA1 A B C GND VCC S
** N=7 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ND3 I3 GND I2 O VCC I1
** N=7 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT XOR2HS I1 I2 O VCC GND
** N=6 EP=5 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MOAI1S B1 B2 GND A1 A2 O VCC
** N=8 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AO112 O C2 C1 VCC B1 GND A1
** N=8 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OR3B2 I1 B1 VCC O B2 GND
** N=7 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AO222 C1 C2 B2 B1 A1 A2 GND VCC O
** N=10 EP=9 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OAI112HS C2 C1 GND B1 O A1 VCC
** N=8 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OR2 I2 I1 VCC GND O
** N=6 EP=5 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OAI12HS B2 B1 GND A1 VCC O
** N=7 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT NR3 I1 VCC I2 I3 O GND
** N=7 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AOI12HS B2 B1 VCC A1 GND O
** N=7 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MAOI1 B1 B2 A1 A2 VCC GND O
** N=8 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OA222 A2 A1 B2 B1 C2 C1 GND VCC O
** N=10 EP=9 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AN2 I1 I2 GND VCC O
** N=6 EP=5 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT XNR2HS I1 I2 O VCC GND
** N=6 EP=5 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_25 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
** N=434 EP=40 IP=2216 FDC=0
X0 53 38 59 39 INV1S $T=460660 800240 0 0 $X=460660 $Y=799860
X1 81 38 55 39 INV1S $T=468720 790160 0 180 $X=467480 $Y=784740
X2 50 38 65 39 INV1S $T=468100 759920 0 0 $X=468100 $Y=759540
X3 64 38 70 39 INV1S $T=475540 770000 1 0 $X=475540 $Y=764580
X4 82 38 100 39 INV1S $T=489800 709520 0 0 $X=489800 $Y=709140
X5 87 38 75 39 INV1S $T=489800 830480 1 0 $X=489800 $Y=825060
X6 83 38 99 39 INV1S $T=492280 729680 1 0 $X=492280 $Y=724260
X7 110 38 102 39 INV1S $T=499720 770000 1 180 $X=498480 $Y=769620
X8 118 38 112 39 INV1S $T=503440 820400 1 180 $X=502200 $Y=820020
X9 53 38 126 39 INV1S $T=507780 790160 1 0 $X=507780 $Y=784740
X10 91 38 117 39 INV1S $T=508400 739760 0 0 $X=508400 $Y=739380
X11 123 38 130 39 INV1S $T=509640 820400 1 0 $X=509640 $Y=814980
X12 149 38 122 39 INV1S $T=516460 770000 0 180 $X=515220 $Y=764580
X13 145 38 150 39 INV1S $T=515220 820400 1 0 $X=515220 $Y=814980
X14 166 38 72 39 INV1S $T=522660 739760 1 180 $X=521420 $Y=739380
X15 131 38 155 39 INV1S $T=521420 810320 1 0 $X=521420 $Y=804900
X16 42 38 172 39 INV1S $T=525140 790160 1 0 $X=525140 $Y=784740
X17 170 38 171 39 INV1S $T=525140 810320 0 0 $X=525140 $Y=809940
X18 146 38 168 39 INV1S $T=525760 719600 0 0 $X=525760 $Y=719220
X19 177 38 132 39 INV1S $T=528240 729680 1 180 $X=527000 $Y=729300
X20 18 38 129 39 INV1S $T=530100 870800 1 180 $X=528860 $Y=870420
X21 49 38 163 39 INV1S $T=533200 719600 1 180 $X=531960 $Y=719220
X22 173 38 195 39 INV1S $T=535680 699440 0 180 $X=534440 $Y=694020
X23 52 38 151 39 INV1S $T=538160 739760 0 0 $X=538160 $Y=739380
X24 47 38 212 39 INV1S $T=540020 790160 0 0 $X=540020 $Y=789780
X25 161 38 135 39 INV1S $T=541260 830480 1 0 $X=541260 $Y=825060
X26 60 38 218 39 INV1S $T=543740 770000 0 0 $X=543740 $Y=769620
X27 45 38 223 39 INV1S $T=547460 800240 1 0 $X=547460 $Y=794820
X28 86 38 232 39 INV1S $T=551180 790160 0 0 $X=551180 $Y=789780
X29 51 38 157 39 INV1S $T=553660 719600 0 0 $X=553660 $Y=719220
X30 168 38 175 39 INV1S $T=556140 749840 1 0 $X=556140 $Y=744420
X31 66 38 247 39 INV1S $T=556140 790160 0 0 $X=556140 $Y=789780
X32 181 38 141 39 INV1S $T=575980 790160 0 0 $X=575980 $Y=789780
X33 196 38 116 39 INV1S $T=581560 770000 1 0 $X=581560 $Y=764580
X34 81 38 288 39 INV1S $T=584660 800240 1 180 $X=583420 $Y=799860
X35 46 38 304 39 INV1S $T=587140 790160 0 0 $X=587140 $Y=789780
X36 73 38 114 39 INV1S $T=594580 810320 0 180 $X=593340 $Y=804900
X37 111 38 106 39 INV1S $T=604500 800240 1 180 $X=603260 $Y=799860
X38 3 38 39 43 BUF1 $T=447640 770000 1 180 $X=445160 $Y=769620
X39 3 38 39 56 BUF1 $T=453840 820400 0 0 $X=453840 $Y=820020
X40 3 38 39 54 BUF1 $T=456320 840560 0 0 $X=456320 $Y=840180
X41 68 38 39 41 BUF1 $T=473680 699440 0 180 $X=471200 $Y=694020
X42 43 38 39 68 BUF1 $T=471200 709520 1 0 $X=471200 $Y=704100
X43 63 38 39 136 BUF1 $T=511500 759920 1 0 $X=511500 $Y=754500
X44 72 38 39 143 BUF1 $T=513360 729680 0 0 $X=513360 $Y=729300
X45 130 38 39 152 BUF1 $T=514600 810320 1 0 $X=514600 $Y=804900
X46 132 38 39 71 BUF1 $T=516460 759920 1 0 $X=516460 $Y=754500
X47 155 38 39 80 BUF1 $T=523280 780080 0 180 $X=520800 $Y=774660
X48 139 38 39 199 BUF1 $T=533820 780080 1 0 $X=533820 $Y=774660
X49 150 38 39 202 BUF1 $T=536300 749840 1 0 $X=536300 $Y=744420
X50 54 38 39 224 BUF1 $T=546840 830480 0 0 $X=546840 $Y=830100
X51 126 38 39 250 BUF1 $T=556140 759920 0 0 $X=556140 $Y=759540
X52 172 38 39 256 BUF1 $T=560480 790160 1 0 $X=560480 $Y=784740
X53 114 38 39 244 BUF1 $T=560480 800240 1 0 $X=560480 $Y=794820
X54 223 38 39 267 BUF1 $T=564820 790160 0 0 $X=564820 $Y=789780
X55 106 38 39 225 BUF1 $T=567920 770000 1 0 $X=567920 $Y=764580
X56 218 38 39 271 BUF1 $T=570400 770000 0 0 $X=570400 $Y=769620
X57 288 38 39 204 BUF1 $T=576600 800240 1 180 $X=574120 $Y=799860
X58 212 38 39 289 BUF1 $T=575980 759920 0 0 $X=575980 $Y=759540
X59 68 38 39 314 BUF1 $T=585900 699440 1 0 $X=585900 $Y=694020
X60 151 38 39 317 BUF1 $T=596440 749840 1 0 $X=596440 $Y=744420
X61 141 38 39 303 BUF1 $T=597060 770000 0 0 $X=597060 $Y=769620
X62 232 38 39 322 BUF1 $T=598300 790160 0 0 $X=598300 $Y=789780
X63 163 38 39 337 BUF1 $T=605740 759920 1 0 $X=605740 $Y=754500
X64 116 38 39 338 BUF1 $T=605740 770000 1 0 $X=605740 $Y=764580
X65 304 38 39 329 BUF1 $T=606360 790160 0 0 $X=606360 $Y=789780
X66 157 38 39 351 BUF1 $T=615040 770000 0 0 $X=615040 $Y=769620
X67 247 38 39 355 BUF1 $T=616280 790160 0 0 $X=616280 $Y=789780
X68 224 38 39 368 BUF1 $T=620000 830480 0 0 $X=620000 $Y=830100
X69 143 38 39 405 BUF1 $T=660920 729680 1 0 $X=660920 $Y=724260
X70 202 38 39 412 BUF1 $T=665880 739760 1 0 $X=665880 $Y=734340
X71 193 38 39 415 BUF1 $T=670220 719600 0 0 $X=670220 $Y=719220
X72 1 2 3 38 39 42 QDFFRBN $T=416020 800240 0 0 $X=416020 $Y=799860
X73 44 2 41 38 39 4 QDFFRBN $T=438340 689360 1 180 $X=426560 $Y=688980
X74 5 2 3 38 39 45 QDFFRBN $T=427180 780080 0 0 $X=427180 $Y=779700
X75 6 2 43 38 39 53 QDFFRBN $T=429040 749840 0 0 $X=429040 $Y=749460
X76 7 2 43 38 39 49 QDFFRBN $T=430280 709520 0 0 $X=430280 $Y=709140
X77 8 2 3 38 39 46 QDFFRBN $T=432140 790160 0 0 $X=432140 $Y=789780
X78 9 2 43 38 39 47 QDFFRBN $T=433380 759920 0 0 $X=433380 $Y=759540
X79 11 2 41 38 39 51 QDFFRBN $T=438340 679280 0 0 $X=438340 $Y=678900
X80 12 2 43 38 39 52 QDFFRBN $T=438960 719600 0 0 $X=438960 $Y=719220
X81 48 2 43 38 39 10 QDFFRBN $T=450740 729680 1 180 $X=438960 $Y=729300
X82 13 2 54 38 39 60 QDFFRBN $T=450740 830480 0 0 $X=450740 $Y=830100
X83 14 2 56 38 39 66 QDFFRBN $T=451360 810320 0 0 $X=451360 $Y=809940
X84 67 2 54 38 39 87 QDFFRBN $T=473060 840560 1 0 $X=473060 $Y=835140
X85 15 2 56 38 39 86 QDFFRBN $T=473680 820400 1 0 $X=473680 $Y=814980
X86 88 2 68 38 39 16 QDFFRBN $T=489180 689360 0 180 $X=477400 $Y=683940
X87 101 2 54 38 39 118 QDFFRBN $T=494140 830480 0 0 $X=494140 $Y=830100
X88 156 2 68 38 39 20 QDFFRBN $T=519560 679280 0 0 $X=519560 $Y=678900
X89 243 2 224 38 39 161 QDFFRBN $T=556760 840560 0 180 $X=544980 $Y=835140
X90 246 2 68 38 39 21 QDFFRBN $T=566060 679280 0 0 $X=566060 $Y=678900
X91 185 2 68 38 39 22 QDFFRBN $T=574740 689360 0 0 $X=574740 $Y=688980
X92 24 2 224 38 39 196 QDFFRBN $T=589620 830480 1 180 $X=577840 $Y=830100
X93 23 2 224 38 39 181 QDFFRBN $T=590240 840560 0 180 $X=578460 $Y=835140
X94 25 2 224 38 39 111 QDFFRBN $T=633020 850640 0 180 $X=621240 $Y=845220
X95 26 2 368 38 39 81 QDFFRBN $T=635500 820400 1 180 $X=623720 $Y=820020
X96 211 2 314 38 39 27 QDFFRBN $T=626820 689360 0 0 $X=626820 $Y=688980
X97 378 2 314 38 39 28 QDFFRBN $T=633020 679280 0 0 $X=633020 $Y=678900
X98 182 2 314 38 39 29 QDFFRBN $T=634260 699440 0 0 $X=634260 $Y=699060
X99 30 2 368 38 39 73 QDFFRBN $T=666500 840560 0 180 $X=654720 $Y=835140
X100 411 2 368 38 39 31 QDFFRBN $T=667120 830480 1 0 $X=667120 $Y=825060
X101 423 2 314 38 39 32 QDFFRBN $T=688200 689360 0 0 $X=688200 $Y=688980
X102 425 2 368 38 39 33 QDFFRBN $T=691300 850640 0 0 $X=691300 $Y=850260
X103 428 2 314 38 39 34 QDFFRBN $T=694400 699440 0 0 $X=694400 $Y=699060
X104 432 2 368 38 39 36 QDFFRBN $T=698120 820400 0 0 $X=698120 $Y=820020
X105 429 2 368 38 39 35 QDFFRBN $T=698740 840560 1 0 $X=698740 $Y=835140
X106 434 2 314 38 39 37 QDFFRBN $T=714860 679280 0 0 $X=714860 $Y=678900
X107 50 63 62 50 39 72 38 AOI22S $T=465000 759920 1 0 $X=465000 $Y=754500
X108 80 71 76 70 39 69 38 AOI22S $T=478640 780080 0 180 $X=474920 $Y=774660
X109 85 63 58 64 39 72 38 AOI22S $T=486080 770000 0 180 $X=482360 $Y=764580
X110 80 71 79 65 39 90 38 AOI22S $T=482980 749840 0 0 $X=482980 $Y=749460
X111 80 71 89 102 39 96 38 AOI22S $T=491040 770000 0 0 $X=491040 $Y=769620
X112 103 63 94 110 39 72 38 AOI22S $T=497860 770000 1 0 $X=497860 $Y=764580
X113 155 132 159 100 39 107 38 AOI22S $T=512740 709520 1 180 $X=509020 $Y=709140
X114 105 136 134 83 39 143 38 AOI22S $T=511500 729680 1 0 $X=511500 $Y=724260
X115 124 136 142 82 39 143 38 AOI22S $T=513360 699440 0 0 $X=513360 $Y=699060
X116 138 136 144 91 39 72 38 AOI22S $T=513360 749840 1 0 $X=513360 $Y=744420
X117 137 136 148 149 39 72 38 AOI22S $T=515220 759920 0 0 $X=515220 $Y=759540
X118 155 132 164 99 39 158 38 AOI22S $T=523900 729680 1 180 $X=520180 $Y=729300
X119 80 71 160 122 39 174 38 AOI22S $T=520800 770000 0 0 $X=520800 $Y=769620
X120 155 132 167 117 39 187 38 AOI22S $T=523900 749840 0 0 $X=523900 $Y=749460
X121 168 175 193 132 39 171 38 AOI22S $T=533200 739760 1 180 $X=529480 $Y=739380
X122 268 290 285 202 39 143 38 AOI22S $T=578460 709520 0 0 $X=578460 $Y=709140
X123 397 376 406 202 39 143 38 AOI22S $T=655960 709520 1 180 $X=652240 $Y=709140
X124 399 407 413 412 39 405 38 AOI22S $T=672700 759920 0 180 $X=668980 $Y=754500
X125 399 394 424 412 39 405 38 AOI22S $T=682000 729680 1 180 $X=678280 $Y=729300
X126 399 421 420 412 39 405 38 AOI22S $T=681380 739760 0 0 $X=681380 $Y=739380
X127 397 427 426 412 39 405 38 AOI22S $T=696260 759920 0 180 $X=692540 $Y=754500
X128 397 431 430 412 39 405 38 AOI22S $T=696880 770000 1 0 $X=696880 $Y=764580
X129 397 422 433 412 39 405 38 AOI22S $T=698740 749840 0 0 $X=698740 $Y=749460
X130 81 77 59 39 38 ND2 $T=480500 800240 1 180 $X=478640 $Y=799860
X131 17 180 129 39 38 ND2 $T=529480 860720 1 180 $X=527620 $Y=860340
X132 240 276 199 39 38 ND2 $T=569780 709520 0 180 $X=567920 $Y=704100
X133 406 434 193 39 38 ND2 $T=667740 709520 1 0 $X=667740 $Y=704100
X134 413 411 415 39 38 ND2 $T=671460 810320 1 0 $X=671460 $Y=804900
X135 424 423 415 39 38 ND2 $T=690060 719600 0 0 $X=690060 $Y=719220
X136 426 429 415 39 38 ND2 $T=695020 810320 1 0 $X=695020 $Y=804900
X137 430 425 415 39 38 ND2 $T=696880 790160 1 0 $X=696880 $Y=784740
X138 420 428 415 39 38 ND2 $T=698120 729680 0 0 $X=698120 $Y=729300
X139 433 432 415 39 38 ND2 $T=699980 800240 0 180 $X=698120 $Y=794820
X140 74 38 47 114 77 39 64 FA1S $T=482980 790160 1 180 $X=471200 $Y=789780
X141 92 38 66 163 93 39 82 FA1S $T=496000 719600 1 180 $X=484220 $Y=719220
X142 93 38 86 151 95 39 83 FA1S $T=496000 739760 0 180 $X=484220 $Y=734340
X143 98 38 45 106 74 39 110 FA1S $T=489180 780080 0 0 $X=489180 $Y=779700
X144 95 38 60 116 109 39 91 FA1S $T=502200 749840 0 180 $X=490420 $Y=744420
X145 109 38 42 141 98 39 149 FA1S $T=504680 780080 1 0 $X=504680 $Y=774660
X146 153 38 73 47 115 39 128 FA1S $T=521420 790160 1 180 $X=509640 $Y=789780
X147 146 38 46 157 92 39 173 FA1S $T=510880 719600 1 0 $X=510880 $Y=714180
X148 184 38 111 45 153 39 190 FA1S $T=525760 800240 1 0 $X=525760 $Y=794820
X149 192 38 181 42 184 39 205 FA1S $T=529480 790160 1 0 $X=529480 $Y=784740
X150 203 38 52 86 198 39 221 FA1S $T=534440 729680 0 0 $X=534440 $Y=729300
X151 198 38 196 60 192 39 217 FA1S $T=535060 759920 0 0 $X=535060 $Y=759540
X152 206 38 49 66 203 39 220 FA1S $T=536300 709520 0 0 $X=536300 $Y=709140
X153 213 38 229 201 219 39 179 FA1S $T=548080 810320 1 180 $X=536300 $Y=809940
X154 226 38 231 214 222 39 200 FA1S $T=554280 749840 0 180 $X=542500 $Y=744420
X155 222 38 236 213 215 39 194 FA1S $T=555520 780080 0 180 $X=543740 $Y=774660
X156 228 38 230 239 226 39 210 FA1S $T=556140 739760 1 180 $X=544360 $Y=739380
X157 230 38 242 255 234 39 214 FA1S $T=556140 759920 0 180 $X=544360 $Y=754500
X158 231 38 241 237 235 39 215 FA1S $T=556140 790160 0 180 $X=544360 $Y=784740
X159 245 38 252 249 228 39 209 FA1S $T=561100 729680 1 180 $X=549320 $Y=729300
X160 240 38 51 46 206 39 238 FA1S $T=550560 709520 1 0 $X=550560 $Y=704100
X161 254 38 258 261 259 39 234 FA1S $T=567920 770000 1 180 $X=556140 $Y=769620
X162 252 38 254 264 251 39 239 FA1S $T=571020 739760 1 180 $X=559240 $Y=739380
X163 262 38 272 301 245 39 248 FA1S $T=571640 719600 1 180 $X=559860 $Y=719220
X164 263 38 265 269 270 39 251 FA1S $T=571640 749840 0 180 $X=559860 $Y=744420
X165 272 38 263 273 274 39 249 FA1S $T=575980 729680 1 180 $X=564200 $Y=729300
X166 277 38 283 281 278 39 264 FA1S $T=578460 780080 0 180 $X=566680 $Y=774660
X167 287 38 275 293 279 39 273 FA1S $T=583420 759920 0 180 $X=571640 $Y=754500
X168 291 38 302 277 286 39 274 FA1S $T=584660 729680 0 180 $X=572880 $Y=724260
X169 298 38 297 294 295 39 286 FA1S $T=580940 780080 1 0 $X=580940 $Y=774660
X170 308 38 316 315 287 39 299 FA1S $T=597680 759920 0 180 $X=585900 $Y=754500
X171 309 38 319 305 311 39 316 FA1S $T=589000 759920 0 0 $X=589000 $Y=759540
X172 310 38 306 320 307 39 315 FA1S $T=589620 790160 1 0 $X=589620 $Y=784740
X173 318 38 291 326 299 39 301 FA1S $T=602640 719600 1 180 $X=590860 $Y=719220
X174 313 38 300 323 298 39 326 FA1S $T=590860 729680 1 0 $X=590860 $Y=724260
X175 328 38 318 334 262 39 290 FA1S $T=608220 709520 1 180 $X=596440 $Y=709140
X176 333 38 339 330 327 39 342 FA1S $T=601400 780080 1 0 $X=601400 $Y=774660
X177 335 38 344 310 309 39 346 FA1S $T=602640 749840 1 0 $X=602640 $Y=744420
X178 345 38 340 336 324 39 332 FA1S $T=617520 739760 1 180 $X=605740 $Y=739380
X179 341 38 342 332 313 39 352 FA1S $T=606360 739760 1 0 $X=606360 $Y=734340
X180 348 38 346 308 352 39 334 FA1S $T=619380 729680 0 180 $X=607600 $Y=724260
X181 347 38 331 350 343 39 356 FA1S $T=609460 800240 1 0 $X=609460 $Y=794820
X182 360 38 353 333 357 39 369 FA1S $T=618140 749840 1 0 $X=618140 $Y=744420
X183 364 38 361 354 362 39 374 FA1S $T=620620 770000 0 0 $X=620620 $Y=769620
X184 366 38 348 359 328 39 376 FA1S $T=621240 719600 0 0 $X=621240 $Y=719220
X185 367 38 374 345 335 39 377 FA1S $T=621860 739760 1 0 $X=621860 $Y=734340
X186 370 38 363 375 358 39 357 FA1S $T=634260 759920 0 180 $X=622480 $Y=754500
X187 372 38 369 341 377 39 359 FA1S $T=635500 729680 0 180 $X=623720 $Y=724260
X188 371 38 379 365 373 39 386 FA1S $T=624960 800240 1 0 $X=624960 $Y=794820
X189 381 38 370 356 360 39 390 FA1S $T=633020 749840 1 0 $X=633020 $Y=744420
X190 389 38 392 367 390 39 382 FA1S $T=649760 739760 1 180 $X=637980 $Y=739380
X191 387 38 380 385 364 39 392 FA1S $T=638600 759920 0 0 $X=638600 $Y=759540
X192 388 38 372 382 366 39 394 FA1S $T=640460 729680 1 0 $X=640460 $Y=724260
X193 391 38 383 347 386 39 393 FA1S $T=641700 800240 1 0 $X=641700 $Y=794820
X194 395 38 387 393 381 39 403 FA1S $T=647900 749840 0 0 $X=647900 $Y=749460
X195 398 38 389 403 388 39 421 FA1S $T=652240 749840 1 0 $X=652240 $Y=744420
X196 408 38 401 404 409 39 417 FA1S $T=662160 780080 1 0 $X=662160 $Y=774660
X197 409 38 384 402 396 39 418 FA1S $T=662780 780080 0 0 $X=662780 $Y=779700
X198 414 38 417 410 416 39 407 FA1S $T=677660 770000 0 180 $X=665880 $Y=764580
X199 410 38 371 418 391 39 419 FA1S $T=665880 790160 0 0 $X=665880 $Y=789780
X200 416 38 419 395 398 39 422 FA1S $T=668980 749840 0 0 $X=668980 $Y=749460
X201 427 38 400 408 414 39 431 FA1S $T=695640 770000 0 0 $X=695640 $Y=769620
X202 140 38 133 17 39 NR2 $T=513360 850640 1 0 $X=513360 $Y=845220
X203 18 38 140 19 39 NR2 $T=513360 860720 0 0 $X=513360 $Y=860340
X204 139 38 176 171 39 NR2 $T=531340 820400 0 180 $X=529480 $Y=814980
X205 204 38 154 126 39 NR2 $T=540640 780080 0 180 $X=538780 $Y=774660
X206 204 38 216 212 39 NR2 $T=541880 800240 1 0 $X=541880 $Y=794820
X207 212 38 227 225 39 NR2 $T=546840 770000 1 0 $X=546840 $Y=764580
X208 126 38 229 106 39 NR2 $T=552420 810320 0 180 $X=550560 $Y=804900
X209 223 38 237 244 39 NR2 $T=554280 800240 1 0 $X=554280 $Y=794820
X210 126 38 208 244 39 NR2 $T=558000 810320 1 0 $X=558000 $Y=804900
X211 126 38 253 141 39 NR2 $T=558620 780080 0 0 $X=558620 $Y=779700
X212 250 38 257 116 39 NR2 $T=559860 749840 0 0 $X=559860 $Y=749460
X213 204 38 241 172 39 NR2 $T=562340 790160 1 180 $X=560480 $Y=789780
X214 204 38 258 218 39 NR2 $T=562340 780080 1 0 $X=562340 $Y=774660
X215 172 38 259 244 39 NR2 $T=564820 790160 1 0 $X=564820 $Y=784740
X216 212 38 260 244 39 NR2 $T=567300 800240 1 180 $X=565440 $Y=799860
X217 267 38 261 225 39 NR2 $T=567920 770000 0 180 $X=566060 $Y=764580
X218 271 38 265 244 39 NR2 $T=571020 790160 0 180 $X=569160 $Y=784740
X219 204 38 284 223 39 NR2 $T=571020 800240 0 180 $X=569160 $Y=794820
X220 218 38 275 225 39 NR2 $T=572260 759920 0 0 $X=572260 $Y=759540
X221 267 38 281 141 39 NR2 $T=573500 790160 1 0 $X=573500 $Y=784740
X222 256 38 278 225 39 NR2 $T=575980 770000 1 180 $X=574120 $Y=769620
X223 250 38 280 163 39 NR2 $T=575980 739760 0 0 $X=575980 $Y=739380
X224 288 38 283 232 39 NR2 $T=578460 790160 1 0 $X=578460 $Y=784740
X225 267 38 294 116 39 NR2 $T=579700 770000 0 0 $X=579700 $Y=769620
X226 232 38 295 114 39 NR2 $T=581560 790160 0 0 $X=581560 $Y=789780
X227 289 38 296 151 39 NR2 $T=582180 739760 0 0 $X=582180 $Y=739380
X228 289 38 266 303 39 NR2 $T=582180 759920 0 0 $X=582180 $Y=759540
X229 288 38 297 247 39 NR2 $T=583420 790160 1 0 $X=583420 $Y=784740
X230 289 38 282 116 39 NR2 $T=584660 749840 1 0 $X=584660 $Y=744420
X231 256 38 293 303 39 NR2 $T=585280 770000 0 0 $X=585280 $Y=769620
X232 288 38 306 304 39 NR2 $T=588380 800240 1 0 $X=588380 $Y=794820
X233 250 38 312 157 39 NR2 $T=589000 739760 0 0 $X=589000 $Y=739380
X234 256 38 305 116 39 NR2 $T=590860 770000 1 180 $X=589000 $Y=769620
X235 250 38 292 151 39 NR2 $T=590240 749840 1 0 $X=590240 $Y=744420
X236 247 38 307 114 39 NR2 $T=592100 790160 0 0 $X=592100 $Y=789780
X237 271 38 311 303 39 NR2 $T=592720 770000 0 0 $X=592720 $Y=769620
X238 267 38 320 317 39 NR2 $T=595820 780080 1 0 $X=595820 $Y=774660
X239 304 38 331 141 39 NR2 $T=595820 800240 1 0 $X=595820 $Y=794820
X240 289 38 321 163 39 NR2 $T=599540 739760 0 0 $X=599540 $Y=739380
X241 157 38 325 289 39 NR2 $T=603260 759920 0 180 $X=601400 $Y=754500
X242 322 38 319 106 39 NR2 $T=602020 770000 1 0 $X=602020 $Y=764580
X243 329 38 327 114 39 NR2 $T=603880 790160 1 180 $X=602020 $Y=789780
X244 256 38 330 317 39 NR2 $T=605120 780080 0 0 $X=605120 $Y=779700
X245 322 38 336 303 39 NR2 $T=608840 759920 0 0 $X=608840 $Y=759540
X246 271 38 339 338 39 NR2 $T=609460 780080 0 0 $X=609460 $Y=779700
X247 355 38 340 106 39 NR2 $T=613180 770000 0 180 $X=611320 $Y=764580
X248 271 38 343 337 39 NR2 $T=611320 790160 0 0 $X=611320 $Y=789780
X249 351 38 350 256 39 NR2 $T=616280 780080 1 180 $X=614420 $Y=779700
X250 267 38 349 337 39 NR2 $T=617520 759920 1 180 $X=615660 $Y=759540
X251 351 38 354 267 39 NR2 $T=618760 780080 0 180 $X=616900 $Y=774660
X252 355 38 358 303 39 NR2 $T=621860 759920 1 180 $X=620000 $Y=759540
X253 256 38 362 337 39 NR2 $T=620000 780080 0 0 $X=620000 $Y=779700
X254 271 38 363 317 39 NR2 $T=624340 759920 0 0 $X=624340 $Y=759540
X255 329 38 361 106 39 NR2 $T=626200 780080 0 180 $X=624340 $Y=774660
X256 351 38 365 271 39 NR2 $T=626200 790160 0 180 $X=624340 $Y=784740
X257 322 38 375 338 39 NR2 $T=629300 759920 0 0 $X=629300 $Y=759540
X258 329 38 379 338 39 NR2 $T=629920 780080 0 0 $X=629920 $Y=779700
X259 322 38 373 337 39 NR2 $T=633640 790160 0 180 $X=631780 $Y=784740
X260 355 38 380 338 39 NR2 $T=637360 770000 0 180 $X=635500 $Y=764580
X261 329 38 384 317 39 NR2 $T=636740 780080 1 0 $X=636740 $Y=774660
X262 355 38 383 317 39 NR2 $T=637360 780080 0 0 $X=637360 $Y=779700
X263 322 38 385 317 39 NR2 $T=644800 770000 0 180 $X=642940 $Y=764580
X264 351 38 402 322 39 NR2 $T=646660 780080 1 180 $X=644800 $Y=779700
X265 329 38 401 337 39 NR2 $T=646040 770000 0 0 $X=646040 $Y=769620
X266 355 38 396 337 39 NR2 $T=649140 790160 0 180 $X=647280 $Y=784740
X267 351 38 404 355 39 NR2 $T=652860 770000 1 0 $X=652860 $Y=764580
X268 351 38 400 329 39 NR2 $T=652860 780080 1 0 $X=652860 $Y=774660
X269 197 38 397 168 39 NR2 $T=654100 719600 0 0 $X=654100 $Y=719220
X270 197 38 399 168 39 NR2 $T=654720 739760 1 0 $X=654720 $Y=734340
X271 70 65 84 39 38 85 HA1 $T=478640 759920 0 0 $X=478640 $Y=759540
X272 102 84 104 39 38 103 HA1 $T=492280 759920 0 0 $X=492280 $Y=759540
X273 99 119 108 39 38 105 HA1 $T=506540 729680 0 180 $X=498480 $Y=724260
X274 100 108 120 39 38 124 HA1 $T=499720 699440 0 0 $X=499720 $Y=699060
X275 117 113 119 39 38 138 HA1 $T=500340 749840 0 0 $X=500340 $Y=749460
X276 122 104 113 39 38 137 HA1 $T=503440 759920 0 0 $X=503440 $Y=759540
X277 195 120 197 39 38 169 HA1 $T=530100 699440 0 0 $X=530100 $Y=699060
X278 208 216 201 39 38 147 HA1 $T=546220 800240 1 180 $X=538160 $Y=799860
X279 227 253 242 39 38 236 HA1 $T=562340 770000 0 180 $X=554280 $Y=764580
X280 266 257 269 39 38 255 HA1 $T=562960 759920 1 0 $X=562960 $Y=754500
X281 282 292 279 39 38 270 HA1 $T=582180 749840 0 180 $X=574120 $Y=744420
X282 284 260 235 39 38 219 HA1 $T=582180 810320 1 180 $X=574120 $Y=809940
X283 296 280 300 39 38 302 HA1 $T=579700 729680 0 0 $X=579700 $Y=729300
X284 321 312 324 39 38 323 HA1 $T=593960 739760 1 0 $X=593960 $Y=734340
X285 349 325 353 39 38 344 HA1 $T=611320 759920 1 0 $X=611320 $Y=754500
X286 118 39 135 123 38 87 ND3 $T=513360 820400 1 180 $X=510880 $Y=820020
X287 118 39 135 145 38 75 ND3 $T=511500 830480 0 0 $X=511500 $Y=830100
X288 118 39 75 162 38 161 ND3 $T=520800 840560 1 0 $X=520800 $Y=835140
X289 161 39 112 131 38 87 ND3 $T=523900 830480 0 180 $X=521420 $Y=825060
X290 19 39 17 178 38 18 ND3 $T=528240 860720 1 0 $X=528240 $Y=855300
X291 87 39 135 170 38 112 ND3 $T=530720 820400 0 0 $X=530720 $Y=820020
X292 161 39 112 177 38 75 ND3 $T=533200 830480 1 180 $X=530720 $Y=830100
X293 285 39 276 378 38 193 ND3 $T=577840 709520 1 0 $X=577840 $Y=704100
X294 47 73 69 38 39 XOR2HS $T=479880 780080 1 180 $X=474300 $Y=779700
X295 53 81 90 38 39 XOR2HS $T=487940 790160 1 0 $X=487940 $Y=784740
X296 66 49 107 38 39 XOR2HS $T=496000 709520 0 0 $X=496000 $Y=709140
X297 45 111 96 38 39 XOR2HS $T=501580 800240 1 180 $X=496000 $Y=799860
X298 86 52 158 38 39 XOR2HS $T=518320 739760 1 0 $X=518320 $Y=734340
X299 46 51 165 38 39 XOR2HS $T=528240 699440 1 180 $X=522660 $Y=699060
X300 42 181 174 38 39 XOR2HS $T=531340 780080 0 180 $X=525760 $Y=774660
X301 60 196 187 38 39 XOR2HS $T=536300 759920 0 180 $X=530720 $Y=754500
X302 197 175 268 38 39 XOR2HS $T=564200 709520 0 0 $X=564200 $Y=709140
X303 78 17 39 78 75 67 38 MOAI1S $T=481740 850640 0 180 $X=478020 $Y=845220
X304 78 18 39 78 112 101 38 MOAI1S $T=497860 850640 0 0 $X=497860 $Y=850260
X305 183 178 39 180 162 78 38 MOAI1S $T=531960 850640 0 180 $X=528240 $Y=845220
X306 78 19 39 78 135 243 38 MOAI1S $T=553040 850640 1 0 $X=553040 $Y=845220
X307 248 202 39 173 177 233 38 MOAI1S $T=557380 719600 0 180 $X=553660 $Y=714180
X308 246 199 238 38 188 39 233 AO112 $T=557380 699440 1 180 $X=552420 $Y=699060
X309 57 58 38 44 76 39 OR3B2 $T=459420 770000 0 0 $X=459420 $Y=769620
X310 61 62 38 48 79 39 OR3B2 $T=464380 749840 1 0 $X=464380 $Y=744420
X311 97 94 38 88 89 39 OR3B2 $T=494140 770000 0 180 $X=490420 $Y=764580
X312 186 148 38 156 160 39 OR3B2 $T=531340 770000 0 180 $X=527620 $Y=764580
X313 191 134 38 182 164 39 OR3B2 $T=533820 729680 0 180 $X=530100 $Y=724260
X314 189 144 38 185 167 39 OR3B2 $T=533820 749840 0 180 $X=530100 $Y=744420
X315 207 142 38 211 159 39 OR3B2 $T=545600 709520 0 180 $X=541880 $Y=704100
X316 128 139 130 111 147 150 39 38 57 AO222 $T=512120 800240 0 0 $X=512120 $Y=799860
X317 90 139 152 73 154 150 39 38 61 AO222 $T=514600 780080 0 0 $X=514600 $Y=779700
X318 155 165 143 169 136 173 39 38 188 AO222 $T=522660 709520 0 0 $X=522660 $Y=709140
X319 190 139 152 181 179 150 39 38 97 AO222 $T=533820 800240 1 180 $X=527620 $Y=799860
X320 205 199 152 196 194 150 39 38 186 AO222 $T=538780 770000 1 180 $X=532580 $Y=769620
X321 217 199 152 52 200 150 39 38 189 AO222 $T=542500 749840 1 180 $X=536300 $Y=749460
X322 220 199 152 51 209 202 39 38 207 AO222 $T=546840 719600 1 180 $X=540640 $Y=719220
X323 221 199 152 49 210 202 39 38 191 AO222 $T=546840 729680 0 180 $X=540640 $Y=724260
X324 177 180 39 121 183 176 38 OAI112HS $T=533820 840560 1 180 $X=529480 $Y=840180
X325 175 162 38 39 166 OR2 $T=527620 749840 0 180 $X=525140 $Y=744420
X326 162 168 39 170 38 63 OAI12HS $T=523280 759920 1 0 $X=523280 $Y=754500
X327 118 38 161 87 139 39 NR3 $T=520180 820400 0 0 $X=520180 $Y=820020
X328 19 18 38 140 39 125 AOI12HS $T=510880 860720 1 0 $X=510880 $Y=855300
X329 17 19 17 129 38 39 127 MAOI1 $T=507160 870800 0 0 $X=507160 $Y=870420
X330 145 133 131 127 123 125 39 38 121 OA222 $T=512740 840560 1 180 $X=507160 $Y=840180
X331 53 81 39 38 115 AN2 $T=499100 790160 1 0 $X=499100 $Y=784740
X332 55 53 50 38 39 XNR2HS $T=460040 780080 1 180 $X=454460 $Y=779700
.ENDS
***************************************
.SUBCKT ICV_26
** N=20 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_27 1 2 3 17 18 44
** N=44 EP=6 IP=10 FDC=0
X0 17 1 3 18 INV1S $T=807240 225680 1 180 $X=806000 $Y=225300
X1 3 1 18 2 BUF1 $T=426560 225680 0 180 $X=424080 $Y=220260
.ENDS
***************************************
.SUBCKT ICV_28 1 8 9 10 11 12 13 36
** N=50 EP=8 IP=16 FDC=0
X0 8 9 9 9 10 11 1 YA2GSD $T=403000 0 0 0 $X=405850 $Y=0
X1 12 11 11 11 13 11 1 YA2GSD $T=511500 0 0 0 $X=514350 $Y=0
.ENDS
***************************************
.SUBCKT ICV_29 1 2 3 4 5 6 9
** N=11 EP=7 IP=12 FDC=0
X0 2 3 3 3 4 XMD $T=231930 1403480 0 180 $X=172160 $Y=1263980
X1 5 1 1 1 6 XMD $T=323740 1403480 0 180 $X=263970 $Y=1263980
.ENDS
***************************************
.SUBCKT INV12CK I O GND VCC
** N=5 EP=4 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_30 2 3 4 5 6 7 9 10
** N=10 EP=8 IP=15 FDC=0
X0 6 9 3 4 BUF1 $T=233120 1173200 1 180 $X=230640 $Y=1172820
X1 7 9 3 6 BUF1 $T=277140 1183280 0 180 $X=274660 $Y=1177860
X2 2 5 3 9 INV12CK $T=220720 1173200 0 0 $X=220720 $Y=1172820
.ENDS
***************************************
.SUBCKT ICV_31 4 5 6 7 8 9 10 11
** N=11 EP=8 IP=15 FDC=0
X0 4 7 10 5 BUF1 $T=228160 941360 0 180 $X=225680 $Y=935940
X1 6 7 10 4 BUF1 $T=228780 1042160 1 180 $X=226300 $Y=1041780
X2 8 9 10 7 INV12CK $T=248620 1082480 0 0 $X=248620 $Y=1082100
.ENDS
***************************************
.SUBCKT ICV_32
** N=7 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_33
** N=6 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_34 4 6 7 8 9 10 12 14
** N=14 EP=8 IP=20 FDC=0
X0 9 6 12 4 BUF1 $T=228160 225680 0 180 $X=225680 $Y=220260
X1 7 6 12 8 BUF1 $T=228160 376880 1 180 $X=225680 $Y=376500
X2 4 6 12 7 BUF1 $T=228780 276080 1 180 $X=226300 $Y=275700
X3 10 6 12 9 BUF1 $T=315580 225680 0 180 $X=313100 $Y=220260
.ENDS
***************************************
.SUBCKT ICV_35 1 2 3 4 5 6 7 8 10
** N=11 EP=9 IP=16 FDC=0
X0 3 4 1 1 5 1 2 YA2GSD $T=186000 0 0 0 $X=188850 $Y=0
X1 6 1 1 7 8 7 2 YA2GSD $T=294500 0 0 0 $X=297350 $Y=0
.ENDS
***************************************
.SUBCKT ICV_36
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_37 1 2 3 4 7
** N=8 EP=5 IP=6 FDC=0
X0 4 3 3 2 1 XMD $T=0 1241270 0 270 $X=0 $Y=1181500
.ENDS
***************************************
.SUBCKT ICV_38 1 2 3 4 5 6 7 8 11
** N=12 EP=9 IP=18 FDC=0
X0 4 5 5 5 1 XMD $T=0 987150 0 270 $X=0 $Y=927380
X1 6 7 5 5 2 XMD $T=0 1071850 0 270 $X=0 $Y=1012080
X2 8 7 7 7 3 XMD $T=0 1156560 0 270 $X=0 $Y=1096790
.ENDS
***************************************
.SUBCKT ICV_39 1 2 3 4 5 8
** N=22 EP=6 IP=12 FDC=0
X0 4 3 3 3 1 XMD $T=0 817750 0 270 $X=0 $Y=757980
X1 5 3 3 3 2 XMD $T=0 902450 0 270 $X=0 $Y=842680
.ENDS
***************************************
.SUBCKT ICV_40 1 2 3 4 5 8
** N=10 EP=6 IP=12 FDC=0
X0 4 2 2 2 1 XMD $T=0 478950 0 270 $X=0 $Y=419180
X1 5 2 2 2 3 XMD $T=0 563650 0 270 $X=0 $Y=503880
.ENDS
***************************************
.SUBCKT ICV_41 1 2 3 4 5 6 7 8 10
** N=12 EP=9 IP=18 FDC=0
X0 4 5 5 5 1 XMD $T=0 224830 0 270 $X=0 $Y=165060
X1 6 7 7 5 2 XMD $T=0 309540 0 270 $X=0 $Y=249770
X2 8 7 7 7 3 XMD $T=0 394250 0 270 $X=0 $Y=334480
.ENDS
***************************************
.SUBCKT ICV_42
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT CHIP data_o[15] data_o[13] data_o[14] data_o[12] data_o[10] data_o[11] data_o[8] data_o[9] data_a_i[3] data_a_i[4] VCC GND data_o[6] data_o[7] data_a_i[0] data_a_i[1] data_a_i[2] data_o[4] data_o[5] inst_i[0]
+ inst_i[1] inst_i[2] data_o[2] data_o[3] clk_p_i reset_n_i data_o[0] data_o[1] data_b_i[7] data_b_i[4] data_b_i[5] data_b_i[6] data_b_i[2] data_b_i[3] data_b_i[0] data_b_i[1] data_a_i[5] data_a_i[6] data_a_i[7]
** N=169 EP=39 IP=529 FDC=0
X1 data_o[15] 95 116 6 169 ICV_2 $T=0 0 0 0 $X=1271600 $Y=1153700
X2 2 3 4 5 6 data_o[13] data_o[14] 169 ICV_3 $T=0 0 0 0 $X=1271600 $Y=927400
X3 9 10 data_o[12] 6 169 ICV_4 $T=0 0 0 0 $X=1271600 $Y=568500
X4 12 13 14 15 6 data_o[10] 120 data_o[11] 169 ICV_5 $T=0 0 0 0 $X=1271600 $Y=391400
X5 18 19 14 20 data_o[8] data_o[9] 121 12 169 ICV_6 $T=0 0 0 0 $X=1271600 $Y=139500
X7 23 data_a_i[3] 96 data_a_i[4] 95 97 169 ICV_8 $T=0 0 0 0 $X=1055400 $Y=1263980
X8 GND 133 23 95 VCC 169 ICV_9 $T=0 0 0 0 $X=1055400 $Y=1153700
X9 VCC 4 95 3 GND 169 ICV_10 $T=0 0 0 0 $X=1055400 $Y=927400
X10 3 9 VCC GND 169 ICV_11 $T=0 0 0 0 $X=1055400 $Y=568500
X11 12 13 14 6 VCC GND 169 ICV_12 $T=0 0 0 0 $X=1055400 $Y=391400
X12 VCC 28 98 37 14 18 20 12 GND 169 ICV_13 $T=0 0 0 0 $X=1055400 $Y=139500
X13 28 14 data_o[6] 98 99 data_o[7] 18 100 169 ICV_14 $T=0 0 0 0 $X=1055400 $Y=-56920
X14 32 33 data_a_i[0] 36 101 data_a_i[1] 102 data_a_i[2] 104 103 169 ICV_15 $T=0 0 0 0 $X=814800 $Y=1263980
X15 GND 36 32 33 133 104 VCC 169 ICV_16 $T=0 0 0 0 $X=814800 $Y=1153700
X17 38 32 VCC GND 169 ICV_18 $T=0 0 0 0 $X=814800 $Y=568500
X19 VCC 38 39 28 GND 169 ICV_20 $T=0 0 0 0 $X=814800 $Y=139500
X20 39 28 data_o[4] 105 37 data_o[5] 106 169 ICV_21 $T=0 0 0 0 $X=814800 $Y=-56920
X21 42 44 36 inst_i[0] 107 inst_i[1] 108 inst_i[2] 109 169 ICV_22 $T=0 0 0 0 $X=355780 $Y=1263980
X22 GND 42 44 36 VCC 169 ICV_23 $T=0 0 0 0 $X=355800 $Y=1153700
X24 59 140 54 117 58 60 65 53 61 64 66 63 55 57 56 118 107 108 109 119
+ 100 105 96 97 103 101 99 19 106 102 2 120 5 15 116 10 121 VCC GND 169
+ ICV_25 $T=0 0 0 0 $X=355800 $Y=568500
X26 VCC 62 122 38 GND 169 ICV_27 $T=0 0 0 0 $X=355800 $Y=139500
X27 37 data_o[2] 62 118 122 data_o[3] 119 169 ICV_28 $T=0 0 0 0 $X=355800 $Y=-56920
X28 42 clk_p_i 78 129 reset_n_i 54 169 ICV_29 $T=0 0 0 0 $X=139500 $Y=1263980
X29 129 GND 77 147 78 42 VCC 169 ICV_30 $T=0 0 0 0 $X=139500 $Y=1153700
X30 130 79 77 VCC 147 140 GND 169 ICV_31 $T=0 0 0 0 $X=139500 $Y=927400
X33 131 VCC 132 80 81 62 GND 169 ICV_34 $T=0 0 0 0 $X=139500 $Y=139500
X34 81 37 data_o[0] 131 64 data_o[1] 62 117 169 ICV_35 $T=0 0 0 0 $X=139500 $Y=-56920
X36 53 77 78 data_b_i[7] 169 ICV_37 $T=0 0 0 0 $X=-56920 $Y=1153700
X37 55 56 57 data_b_i[4] 130 data_b_i[5] 77 data_b_i[6] 169 ICV_38 $T=0 0 0 0 $X=-56920 $Y=927380
X38 58 59 79 data_b_i[2] data_b_i[3] 169 ICV_39 $T=0 0 0 0 $X=-56920 $Y=568500
X39 60 80 61 data_b_i[0] data_b_i[1] 169 ICV_40 $T=0 0 0 0 $X=-56920 $Y=391400
X40 63 65 66 data_a_i[5] 131 data_a_i[6] 132 data_a_i[7] 169 ICV_41 $T=0 0 0 0 $X=-56920 $Y=139500
.ENDS
***************************************
