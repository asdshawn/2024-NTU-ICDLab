* SPICE NETLIST
***************************************

.SUBCKT L POS NEG SUB
.ENDS
***************************************
.SUBCKT YA2GSD O E2 E8 E4 I SR E
** N=8 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_1 1 2 3 4 5
** N=5 EP=5 IP=8 FDC=0
X0 1 2 2 2 3 2 4 YA2GSD $T=0 0 0 0 $X=2850 $Y=0
.ENDS
***************************************
.SUBCKT ICV_2
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_3 1 2 3 4 5
** N=6 EP=5 IP=8 FDC=0
X0 1 2 2 2 3 2 4 YA2GSD $T=1349740 1096780 0 90 $X=1210240 $Y=1099630
.ENDS
***************************************
.SUBCKT ICV_4 1 2 3 4 7
** N=8 EP=5 IP=8 FDC=0
X0 3 1 1 1 2 1 4 YA2GSD $T=1349740 983520 0 90 $X=1210240 $Y=986370
.ENDS
***************************************
.SUBCKT ICV_5 1 2 4 5 9
** N=10 EP=5 IP=8 FDC=0
X0 4 1 1 1 5 1 2 YA2GSD $T=1349740 757020 0 90 $X=1210240 $Y=759870
.ENDS
***************************************
.SUBCKT ICV_6
** N=13 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_7 2 3 4 5 11
** N=12 EP=5 IP=8 FDC=0
X0 2 3 3 3 4 3 5 YA2GSD $T=1349740 417270 0 90 $X=1210240 $Y=420120
.ENDS
***************************************
.SUBCKT ICV_8 1 2 3 4 5 6 7 8
** N=10 EP=8 IP=16 FDC=0
X0 2 3 3 3 1 3 4 YA2GSD $T=1349740 190760 0 90 $X=1210240 $Y=193610
X1 5 6 6 6 7 6 4 YA2GSD $T=1349740 304020 0 90 $X=1210240 $Y=306870
.ENDS
***************************************
.SUBCKT ICV_9
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT XMD I SMT PU PD O
** N=6 EP=5 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_10 1 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26
+ 47
** N=66 EP=21 IP=46 FDC=0
X0 11 10 9 9 12 9 13 YA2GSD $T=1045810 1350160 0 180 $X=986040 $Y=1210660
X1 14 10 10 10 15 10 13 YA2GSD $T=1159020 1350160 0 180 $X=1099250 $Y=1210660
X2 16 17 17 17 18 XMD $T=253340 1350160 0 180 $X=193570 $Y=1210660
X3 19 1 1 1 20 XMD $T=366550 1350160 0 180 $X=306780 $Y=1210660
X4 21 8 1 1 22 XMD $T=706180 1350160 0 180 $X=646410 $Y=1210660
X5 23 8 8 8 24 XMD $T=819390 1350160 0 180 $X=759620 $Y=1210660
X6 25 9 9 8 26 XMD $T=932600 1350160 0 180 $X=872830 $Y=1210660
.ENDS
***************************************
.SUBCKT TIE0 O VCC GND
** N=4 EP=3 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT BUF1S I GND VCC O
** N=5 EP=4 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT BUF1 I VCC GND O
** N=5 EP=4 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT QDFFRBN D CK RB VCC GND Q
** N=7 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT INV1S I VCC O GND
** N=5 EP=4 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MXL2HS B S OB A VCC GND
** N=7 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT INV8 O I GND VCC
** N=5 EP=4 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT INV12CK I O GND VCC
** N=5 EP=4 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_11 1 2 3 5 6 7 8 9 10 14 15 16 17 21 22 23 24 25 26 27
+ 28 29 30 31 32 33 34 35 36 37 38 39 40 41 42 43 44 45 46 47
+ 48 49 50 51 52 53 54 55 56 83
** N=111 EP=50 IP=296 FDC=0
X0 56 3 2 TIE0 $T=1129640 1112280 1 180 $X=1127780 $Y=1111900
X1 1 2 3 7 BUF1S $T=226300 1122360 0 180 $X=223820 $Y=1116940
X2 8 2 3 1 BUF1S $T=325500 1122360 1 180 $X=323020 $Y=1121980
X3 54 2 3 38 BUF1S $T=904580 1122360 1 180 $X=902100 $Y=1121980
X4 56 2 3 55 BUF1S $T=1129020 1122360 1 180 $X=1126540 $Y=1121980
X5 31 3 2 85 BUF1 $T=646040 1082040 0 180 $X=643560 $Y=1076620
X6 38 3 2 8 BUF1 $T=679520 1122360 1 180 $X=677040 $Y=1121980
X7 55 3 2 54 BUF1 $T=1029820 1122360 1 180 $X=1027340 $Y=1121980
X8 17 16 15 3 2 14 QDFFRBN $T=517080 1082040 0 180 $X=505300 $Y=1076620
X9 89 29 27 3 2 87 QDFFRBN $T=633020 1092120 0 180 $X=621240 $Y=1086700
X10 91 29 27 3 2 93 QDFFRBN $T=634260 1092120 1 0 $X=634260 $Y=1086700
X11 94 29 27 3 2 96 QDFFRBN $T=646660 1092120 1 0 $X=646660 $Y=1086700
X12 97 33 35 3 2 98 QDFFRBN $T=659680 1082040 0 0 $X=659680 $Y=1081660
X13 34 33 35 3 2 36 QDFFRBN $T=661540 1082040 1 0 $X=661540 $Y=1076620
X14 99 33 35 3 2 100 QDFFRBN $T=672080 1082040 0 0 $X=672080 $Y=1081660
X15 102 33 35 3 2 104 QDFFRBN $T=685100 1082040 0 0 $X=685100 $Y=1081660
X16 107 33 43 3 2 105 QDFFRBN $T=711140 1082040 1 180 $X=699360 $Y=1081660
X17 110 33 43 3 2 108 QDFFRBN $T=725400 1082040 0 180 $X=713620 $Y=1076620
X18 46 33 43 3 2 44 QDFFRBN $T=738420 1082040 0 180 $X=726640 $Y=1076620
X19 47 33 48 3 2 49 QDFFRBN $T=738420 1082040 1 0 $X=738420 $Y=1076620
X20 51 50 48 3 2 111 QDFFRBN $T=761980 1082040 0 180 $X=750200 $Y=1076620
X21 52 50 48 3 2 53 QDFFRBN $T=763220 1082040 1 0 $X=763220 $Y=1076620
X22 24 3 23 2 INV1S $T=610080 1082040 1 0 $X=610080 $Y=1076620
X23 25 3 84 2 INV1S $T=613800 1082040 1 0 $X=613800 $Y=1076620
X24 87 3 88 2 INV1S $T=626820 1082040 0 0 $X=626820 $Y=1081660
X25 30 3 86 2 INV1S $T=631160 1082040 0 180 $X=629920 $Y=1076620
X26 93 3 90 2 INV1S $T=644800 1082040 1 180 $X=643560 $Y=1081660
X27 96 3 92 2 INV1S $T=652860 1082040 1 180 $X=651620 $Y=1081660
X28 98 3 95 2 INV1S $T=657200 1082040 1 180 $X=655960 $Y=1081660
X29 100 3 37 2 INV1S $T=676420 1082040 0 180 $X=675180 $Y=1076620
X30 40 3 103 2 INV1S $T=690680 1082040 1 0 $X=690680 $Y=1076620
X31 104 3 101 2 INV1S $T=695020 1082040 0 180 $X=693780 $Y=1076620
X32 105 3 106 2 INV1S $T=706180 1082040 1 0 $X=706180 $Y=1076620
X33 108 3 109 2 INV1S $T=719200 1082040 0 0 $X=719200 $Y=1081660
X34 111 3 45 2 INV1S $T=750200 1082040 0 0 $X=750200 $Y=1081660
X35 23 22 21 84 3 2 MXL2HS $T=606980 1082040 0 180 $X=601400 $Y=1076620
X36 84 85 26 86 3 2 MXL2HS $T=616280 1082040 1 0 $X=616280 $Y=1076620
X37 86 85 28 88 3 2 MXL2HS $T=623100 1082040 1 0 $X=623100 $Y=1076620
X38 88 85 89 90 3 2 MXL2HS $T=629920 1082040 0 0 $X=629920 $Y=1081660
X39 90 85 91 92 3 2 MXL2HS $T=636740 1082040 0 0 $X=636740 $Y=1081660
X40 92 31 94 95 3 2 MXL2HS $T=647280 1082040 1 0 $X=647280 $Y=1076620
X41 95 31 97 32 3 2 MXL2HS $T=654100 1082040 1 0 $X=654100 $Y=1076620
X42 37 39 99 101 3 2 MXL2HS $T=677660 1082040 1 0 $X=677660 $Y=1076620
X43 101 39 102 103 3 2 MXL2HS $T=683860 1082040 1 0 $X=683860 $Y=1076620
X44 103 41 42 106 3 2 MXL2HS $T=697500 1082040 1 0 $X=697500 $Y=1076620
X45 106 41 107 109 3 2 MXL2HS $T=713000 1082040 0 0 $X=713000 $Y=1081660
X46 109 41 110 45 3 2 MXL2HS $T=722300 1082040 0 0 $X=722300 $Y=1081660
X47 10 9 2 3 INV8 $T=333560 1112280 1 180 $X=327360 $Y=1111900
X48 5 6 2 3 INV12CK $T=220100 1122360 0 0 $X=220100 $Y=1121980
.ENDS
***************************************
.SUBCKT AN2 I1 I2 GND VCC O
** N=6 EP=5 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ND2 I1 O I2 GND VCC
** N=6 EP=5 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OAI12HS B2 B1 GND A1 VCC O
** N=7 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT NR2T O I2 GND I1 VCC
** N=6 EP=5 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ND3 I3 GND I2 O VCC I1
** N=7 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT XNR2HS I1 I2 O VCC GND
** N=6 EP=5 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT XOR2H I1 I2 O GND VCC
** N=6 EP=5 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT NR2 I1 VCC O I2 GND
** N=6 EP=5 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT NR2P I1 VCC I2 GND O
** N=6 EP=5 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MOAI1 B1 B2 GND A1 O A2 VCC
** N=8 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ND2P I2 GND I1 O VCC
** N=6 EP=5 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MAO222 B1 A1 C1 GND VCC O
** N=7 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT FA1 S B VCC A CI GND CO
** N=8 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OR2 I2 I1 VCC GND O
** N=6 EP=5 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AOI12HS B2 B1 VCC A1 GND O
** N=7 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT XOR2HS I1 I2 O VCC GND
** N=6 EP=5 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MOAI1S B1 B2 GND A1 A2 O VCC
** N=8 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ND2S I1 O I2 VCC GND
** N=6 EP=5 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MOAI1H B1 B2 GND A1 O A2 VCC
** N=8 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT INV2 I O GND VCC
** N=5 EP=4 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT BUF2 I O GND VCC
** N=5 EP=4 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AO22 O A2 A1 VCC B1 B2 GND
** N=8 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT INV3 I O GND VCC
** N=5 EP=4 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT BUF6 I O GND VCC
** N=5 EP=4 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OAI22S B2 GND B1 A2 O A1 VCC
** N=8 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT FA1S CO VCC A B CI GND S
** N=8 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT INV4 I O GND VCC
** N=5 EP=4 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT NR3HP O I3 I2 I1 GND VCC
** N=7 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OR2T I2 I1 GND O VCC
** N=6 EP=5 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AOI13HS B3 O B2 B1 VCC A1 GND
** N=8 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT NR3 I1 VCC I2 I3 O GND
** N=7 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OA12 B2 B1 A1 GND VCC O
** N=7 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OAI22H B2 B1 GND A2 O A1 VCC
** N=8 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OAI112H C2 C1 GND B1 O A1 VCC
** N=8 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT QDFFRBP D CK RB Q GND VCC
** N=7 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT QDFFRBS D CK RB VCC GND Q
** N=7 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OAI222S C1 C2 GND B1 B2 VCC A1 O A2
** N=10 EP=9 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_12 1 2 3 4 5 6 7 8 9 10 11
** N=11 EP=11 IP=14 FDC=0
X0 1 2 3 4 5 6 QDFFRBN $T=0 0 0 0 $X=0 $Y=-380
X1 7 8 9 4 5 10 QDFFRBN $T=11780 0 0 0 $X=11780 $Y=-380
.ENDS
***************************************
.SUBCKT BUF3 I VCC GND O
** N=5 EP=4 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT INV6 I O GND VCC
** N=5 EP=4 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_13 1 2 3 4 5 6 7 8 9
** N=9 EP=9 IP=12 FDC=0
X0 1 2 3 4 5 6 QDFFRBN $T=0 0 0 0 $X=0 $Y=-380
X1 7 4 8 5 INV1S $T=12400 0 0 0 $X=12400 $Y=-380
.ENDS
***************************************
.SUBCKT ICV_14 1 2 3 4 5 6 7 8 9 10 11
** N=11 EP=11 IP=14 FDC=0
X0 1 2 3 4 5 6 QDFFRBN $T=0 0 0 0 $X=0 $Y=-380
X1 7 8 9 4 5 10 QDFFRBN $T=12400 0 0 0 $X=12400 $Y=-380
.ENDS
***************************************
.SUBCKT BUF4CK I GND O VCC
** N=5 EP=4 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_15 1 2 3 4 5 6 7 8 9
** N=9 EP=9 IP=12 FDC=0
X0 3 2 4 1 INV1S $T=0 0 0 0 $X=0 $Y=-380
X1 5 6 7 8 2 1 MXL2HS $T=-6200 0 0 0 $X=-6200 $Y=-380
.ENDS
***************************************
.SUBCKT INV8CK I O GND VCC
** N=5 EP=4 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT BUF4 I O GND VCC
** N=5 EP=4 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT INV4CK I O GND VCC
** N=5 EP=4 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_16 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140
+ 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160
+ 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180
+ 181 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200
+ 201 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220
+ 221 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240
+ 241 242 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 259 260
+ 261 262 263 264 265 266 267 268 269 270 271 272 273 274 275 276 277 278 279 280
+ 281 282 293
** N=2314 EP=283 IP=13117 FDC=0
X0 1908 1 2 1963 BUF1S $T=789260 910680 1 180 $X=786780 $Y=910300
X1 1908 1 2 2007 BUF1S $T=792360 910680 0 0 $X=792360 $Y=910300
X2 280 1 2 281 BUF1S $T=1127160 900600 0 0 $X=1127160 $Y=900220
X3 282 1 2 280 BUF1S $T=1129640 1011480 1 180 $X=1127160 $Y=1011100
X4 4 2 1 3 BUF1 $T=224440 991320 1 180 $X=221960 $Y=990940
X5 5 2 1 323 BUF1 $T=374480 920760 1 0 $X=374480 $Y=915340
X6 303 2 1 5 BUF1 $T=377580 930840 0 180 $X=375100 $Y=925420
X7 11 2 1 308 BUF1 $T=378200 910680 0 180 $X=375720 $Y=905260
X8 324 2 1 303 BUF1 $T=378200 951000 1 180 $X=375720 $Y=950620
X9 329 2 1 318 BUF1 $T=381920 951000 1 180 $X=379440 $Y=950620
X10 324 2 1 335 BUF1 $T=380060 981240 0 0 $X=380060 $Y=980860
X11 335 2 1 356 BUF1 $T=386260 961080 1 0 $X=386260 $Y=955660
X12 329 2 1 305 BUF1 $T=386880 940920 0 0 $X=386880 $Y=940540
X13 323 2 1 378 BUF1 $T=395560 920760 1 0 $X=395560 $Y=915340
X14 370 2 1 329 BUF1 $T=399280 951000 0 0 $X=399280 $Y=950620
X15 323 2 1 21 BUF1 $T=401760 910680 0 0 $X=401760 $Y=910300
X16 343 2 1 372 BUF1 $T=405480 981240 1 0 $X=405480 $Y=975820
X17 370 2 1 373 BUF1 $T=412920 971160 0 180 $X=410440 $Y=965740
X18 373 2 1 358 BUF1 $T=413540 991320 0 180 $X=411060 $Y=985900
X19 373 2 1 440 BUF1 $T=414780 981240 1 0 $X=414780 $Y=975820
X20 452 2 1 370 BUF1 $T=420980 951000 1 180 $X=418500 $Y=950620
X21 23 2 1 428 BUF1 $T=420360 910680 1 0 $X=420360 $Y=905260
X22 361 2 1 460 BUF1 $T=420360 1001400 1 0 $X=420360 $Y=995980
X23 25 2 1 23 BUF1 $T=425940 900600 1 180 $X=423460 $Y=900220
X24 356 2 1 453 BUF1 $T=424700 951000 0 0 $X=424700 $Y=950620
X25 475 2 1 418 BUF1 $T=427800 1031640 0 180 $X=425320 $Y=1026220
X26 453 2 1 470 BUF1 $T=434000 930840 0 0 $X=434000 $Y=930460
X27 510 2 1 361 BUF1 $T=437100 1011480 0 180 $X=434620 $Y=1006060
X28 407 2 1 510 BUF1 $T=436480 1021560 0 0 $X=436480 $Y=1021180
X29 25 2 1 521 BUF1 $T=437100 900600 0 0 $X=437100 $Y=900220
X30 452 2 1 519 BUF1 $T=438340 951000 0 0 $X=438340 $Y=950620
X31 343 2 1 525 BUF1 $T=438340 971160 1 0 $X=438340 $Y=965740
X32 510 2 1 523 BUF1 $T=438340 1011480 1 0 $X=438340 $Y=1006060
X33 475 2 1 481 BUF1 $T=438960 1031640 1 0 $X=438960 $Y=1026220
X34 401 2 1 520 BUF1 $T=440200 1041720 1 0 $X=440200 $Y=1036300
X35 560 2 1 452 BUF1 $T=448260 940920 0 180 $X=445780 $Y=935500
X36 525 2 1 563 BUF1 $T=447020 961080 0 0 $X=447020 $Y=960700
X37 520 2 1 576 BUF1 $T=449500 1041720 1 0 $X=449500 $Y=1036300
X38 560 2 1 550 BUF1 $T=453840 920760 1 180 $X=451360 $Y=920380
X39 578 2 1 466 BUF1 $T=455700 1001400 0 180 $X=453220 $Y=995980
X40 520 2 1 601 BUF1 $T=455700 1061880 0 0 $X=455700 $Y=1061500
X41 591 2 1 475 BUF1 $T=458800 1011480 1 180 $X=456320 $Y=1011100
X42 37 2 1 34 BUF1 $T=459420 910680 0 180 $X=456940 $Y=905260
X43 525 2 1 622 BUF1 $T=463140 940920 0 0 $X=463140 $Y=940540
X44 591 2 1 578 BUF1 $T=463760 1011480 1 0 $X=463760 $Y=1006060
X45 591 2 1 605 BUF1 $T=463760 1031640 1 0 $X=463760 $Y=1026220
X46 661 2 1 597 BUF1 $T=474920 930840 1 180 $X=472440 $Y=930460
X47 661 2 1 37 BUF1 $T=473060 910680 1 0 $X=473060 $Y=905260
X48 622 2 1 672 BUF1 $T=477400 951000 0 180 $X=474920 $Y=945580
X49 675 2 1 591 BUF1 $T=474920 1011480 1 0 $X=474920 $Y=1006060
X50 605 2 1 686 BUF1 $T=476780 1041720 1 0 $X=476780 $Y=1036300
X51 696 2 1 643 BUF1 $T=482360 1041720 0 180 $X=479880 $Y=1036300
X52 661 2 1 704 BUF1 $T=481120 910680 1 0 $X=481120 $Y=905260
X53 622 2 1 661 BUF1 $T=481120 930840 1 0 $X=481120 $Y=925420
X54 694 2 1 585 BUF1 $T=484220 1001400 0 180 $X=481740 $Y=995980
X55 672 2 1 702 BUF1 $T=485460 961080 1 0 $X=485460 $Y=955660
X56 694 2 1 733 BUF1 $T=489180 1001400 1 0 $X=489180 $Y=995980
X57 696 2 1 750 BUF1 $T=490420 1041720 1 0 $X=490420 $Y=1036300
X58 696 2 1 746 BUF1 $T=491040 1011480 0 0 $X=491040 $Y=1011100
X59 601 2 1 42 BUF1 $T=491040 1061880 0 0 $X=491040 $Y=1061500
X60 753 2 1 715 BUF1 $T=496000 920760 1 180 $X=493520 $Y=920380
X61 715 2 1 650 BUF1 $T=496620 940920 0 180 $X=494140 $Y=935500
X62 704 2 1 47 BUF1 $T=500960 910680 0 180 $X=498480 $Y=905260
X63 53 2 1 675 BUF1 $T=512740 1001400 1 180 $X=510260 $Y=1001020
X64 53 2 1 753 BUF1 $T=513360 930840 0 180 $X=510880 $Y=925420
X65 53 2 1 560 BUF1 $T=512740 930840 0 0 $X=512740 $Y=930460
X66 560 2 1 840 BUF1 $T=515220 930840 1 0 $X=515220 $Y=925420
X67 900 2 1 797 BUF1 $T=526380 1031640 0 180 $X=523900 $Y=1026220
X68 59 2 1 856 BUF1 $T=532580 900600 1 180 $X=530100 $Y=900220
X69 912 2 1 900 BUF1 $T=533820 1031640 0 180 $X=531340 $Y=1026220
X70 367 2 1 891 BUF1 $T=533200 1071960 0 0 $X=533200 $Y=1071580
X71 917 2 1 59 BUF1 $T=536920 900600 1 180 $X=534440 $Y=900220
X72 874 2 1 931 BUF1 $T=535060 940920 1 0 $X=535060 $Y=935500
X73 840 2 1 924 BUF1 $T=545600 930840 0 0 $X=545600 $Y=930460
X74 862 2 1 1007 BUF1 $T=553660 1001400 0 0 $X=553660 $Y=1001020
X75 924 2 1 997 BUF1 $T=558000 930840 0 0 $X=558000 $Y=930460
X76 931 2 1 967 BUF1 $T=561100 940920 0 180 $X=558620 $Y=935500
X77 955 2 1 1013 BUF1 $T=562340 1041720 1 0 $X=562340 $Y=1036300
X78 1027 2 1 1061 BUF1 $T=566060 961080 0 0 $X=566060 $Y=960700
X79 1007 2 1 1077 BUF1 $T=568540 1021560 0 0 $X=568540 $Y=1021180
X80 1027 2 1 1084 BUF1 $T=573500 991320 0 0 $X=573500 $Y=990940
X81 1128 2 1 1042 BUF1 $T=586520 971160 1 180 $X=584040 $Y=970780
X82 1084 2 1 1142 BUF1 $T=585900 1011480 0 0 $X=585900 $Y=1011100
X83 1084 2 1 1149 BUF1 $T=586520 1001400 0 0 $X=586520 $Y=1001020
X84 1128 2 1 1152 BUF1 $T=589000 971160 1 0 $X=589000 $Y=965740
X85 1045 2 1 71 BUF1 $T=590860 900600 0 0 $X=590860 $Y=900220
X86 1152 2 1 1175 BUF1 $T=593960 971160 1 0 $X=593960 $Y=965740
X87 1069 2 1 1187 BUF1 $T=595200 1051800 1 0 $X=595200 $Y=1046380
X88 68 2 1 1193 BUF1 $T=597680 900600 0 0 $X=597680 $Y=900220
X89 1152 2 1 1222 BUF1 $T=602020 991320 1 0 $X=602020 $Y=985900
X90 1222 2 1 1162 BUF1 $T=608220 1001400 0 180 $X=605740 $Y=995980
X91 1175 2 1 1279 BUF1 $T=621860 961080 0 0 $X=621860 $Y=960700
X92 1222 2 1 1288 BUF1 $T=622480 1011480 1 0 $X=622480 $Y=1006060
X93 1300 2 1 1259 BUF1 $T=624960 910680 1 0 $X=624960 $Y=905260
X94 1237 2 1 1217 BUF1 $T=624960 981240 0 0 $X=624960 $Y=980860
X95 1187 2 1 1235 BUF1 $T=626820 1041720 1 0 $X=626820 $Y=1036300
X96 1217 2 1 1321 BUF1 $T=628680 961080 0 0 $X=628680 $Y=960700
X97 91 2 1 1213 BUF1 $T=631780 1071960 0 180 $X=629300 $Y=1066540
X98 1237 2 1 1296 BUF1 $T=629920 991320 1 0 $X=629920 $Y=985900
X99 1279 2 1 1298 BUF1 $T=631160 961080 0 0 $X=631160 $Y=960700
X100 1288 2 1 1188 BUF1 $T=634880 1011480 1 180 $X=632400 $Y=1011100
X101 1187 2 1 1340 BUF1 $T=633640 1051800 0 0 $X=633640 $Y=1051420
X102 94 2 1 1300 BUF1 $T=637980 900600 1 180 $X=635500 $Y=900220
X103 1296 2 1 1350 BUF1 $T=637360 991320 1 0 $X=637360 $Y=985900
X104 90 2 1 1361 BUF1 $T=638600 920760 1 0 $X=638600 $Y=915340
X105 1288 2 1 1372 BUF1 $T=641080 1021560 1 0 $X=641080 $Y=1016140
X106 1288 2 1 1351 BUF1 $T=642940 1011480 1 0 $X=642940 $Y=1006060
X107 1345 2 1 94 BUF1 $T=645420 920760 1 0 $X=645420 $Y=915340
X108 1322 2 1 97 BUF1 $T=647280 1061880 0 0 $X=647280 $Y=1061500
X109 1340 2 1 1384 BUF1 $T=647900 1051800 0 0 $X=647900 $Y=1051420
X110 1340 2 1 1417 BUF1 $T=651000 1061880 0 0 $X=651000 $Y=1061500
X111 97 2 1 1428 BUF1 $T=654100 1071960 1 0 $X=654100 $Y=1066540
X112 1344 2 1 1434 BUF1 $T=658440 1021560 0 0 $X=658440 $Y=1021180
X113 1428 2 1 1424 BUF1 $T=658440 1061880 1 0 $X=658440 $Y=1056460
X114 1420 2 1 1403 BUF1 $T=665260 971160 0 180 $X=662780 $Y=965740
X115 1424 2 1 1471 BUF1 $T=664640 1031640 1 0 $X=664640 $Y=1026220
X116 1420 2 1 1477 BUF1 $T=666500 971160 1 0 $X=666500 $Y=965740
X117 1434 2 1 1454 BUF1 $T=667740 1011480 1 0 $X=667740 $Y=1006060
X118 1420 2 1 1456 BUF1 $T=670840 940920 0 0 $X=670840 $Y=940540
X119 124 2 1 1441 BUF1 $T=682620 910680 0 180 $X=680140 $Y=905260
X120 1477 2 1 1515 BUF1 $T=681380 971160 0 0 $X=681380 $Y=970780
X121 1428 2 1 1534 BUF1 $T=683240 1061880 1 0 $X=683240 $Y=1056460
X122 1534 2 1 120 BUF1 $T=685720 1071960 1 0 $X=685720 $Y=1066540
X123 124 2 1 1567 BUF1 $T=687580 910680 0 0 $X=687580 $Y=910300
X124 1581 2 1 1486 BUF1 $T=693160 981240 1 180 $X=690680 $Y=980860
X125 1534 2 1 1556 BUF1 $T=690680 1051800 0 0 $X=690680 $Y=1051420
X126 1534 2 1 1553 BUF1 $T=691920 1041720 1 0 $X=691920 $Y=1036300
X127 1513 2 1 1581 BUF1 $T=696260 981240 0 0 $X=696260 $Y=980860
X128 1585 2 1 1617 BUF1 $T=703700 940920 0 0 $X=703700 $Y=940540
X129 1635 2 1 1602 BUF1 $T=704320 961080 1 0 $X=704320 $Y=955660
X130 1477 2 1 1635 BUF1 $T=708660 971160 1 180 $X=706180 $Y=970780
X131 1578 2 1 1625 BUF1 $T=706800 1061880 0 0 $X=706800 $Y=1061500
X132 1657 2 1 1503 BUF1 $T=709900 1001400 1 180 $X=707420 $Y=1001020
X133 1553 2 1 1649 BUF1 $T=708660 1031640 0 0 $X=708660 $Y=1031260
X134 1657 2 1 1621 BUF1 $T=712380 991320 0 180 $X=709900 $Y=985900
X135 1556 2 1 129 BUF1 $T=709900 1071960 1 0 $X=709900 $Y=1066540
X136 1625 2 1 130 BUF1 $T=711140 1061880 0 0 $X=711140 $Y=1061500
X137 1635 2 1 1657 BUF1 $T=717960 981240 1 180 $X=715480 $Y=980860
X138 1657 2 1 1702 BUF1 $T=716100 1001400 0 0 $X=716100 $Y=1001020
X139 1635 2 1 1693 BUF1 $T=717340 971160 1 0 $X=717340 $Y=965740
X140 1691 2 1 1624 BUF1 $T=719820 1041720 1 180 $X=717340 $Y=1041340
X141 1617 2 1 1603 BUF1 $T=720440 930840 1 180 $X=717960 $Y=930460
X142 1617 2 1 1703 BUF1 $T=718580 920760 0 0 $X=718580 $Y=920380
X143 1756 2 1 1738 BUF1 $T=732840 1061880 0 180 $X=730360 $Y=1056460
X144 1666 2 1 1685 BUF1 $T=732220 971160 0 0 $X=732220 $Y=970780
X145 1734 2 1 1691 BUF1 $T=734700 1041720 1 180 $X=732220 $Y=1041340
X146 1685 2 1 1732 BUF1 $T=732840 991320 1 0 $X=732840 $Y=985900
X147 1322 2 1 1782 BUF1 $T=738420 991320 1 0 $X=738420 $Y=985900
X148 1734 2 1 1744 BUF1 $T=738420 1031640 1 0 $X=738420 $Y=1026220
X149 1736 2 1 1759 BUF1 $T=741520 951000 1 180 $X=739040 $Y=950620
X150 1703 2 1 156 BUF1 $T=744000 900600 1 180 $X=741520 $Y=900220
X151 1703 2 1 1785 BUF1 $T=743380 910680 0 0 $X=743380 $Y=910300
X152 1703 2 1 157 BUF1 $T=744000 900600 0 0 $X=744000 $Y=900220
X153 157 2 1 160 BUF1 $T=747720 900600 0 0 $X=747720 $Y=900220
X154 1744 2 1 1806 BUF1 $T=748960 1021560 0 0 $X=748960 $Y=1021180
X155 1756 2 1 164 BUF1 $T=752060 1071960 1 0 $X=752060 $Y=1066540
X156 1782 2 1 1857 BUF1 $T=756400 1021560 1 0 $X=756400 $Y=1016140
X157 1857 2 1 1771 BUF1 $T=760120 1041720 0 180 $X=757640 $Y=1036300
X158 1808 2 1 1769 BUF1 $T=758880 930840 0 0 $X=758880 $Y=930460
X159 1871 2 1 1803 BUF1 $T=763840 961080 1 180 $X=761360 $Y=960700
X160 1808 2 1 1864 BUF1 $T=761980 920760 1 0 $X=761980 $Y=915340
X161 1865 2 1 1773 BUF1 $T=764460 1061880 1 180 $X=761980 $Y=1061500
X162 1857 2 1 1899 BUF1 $T=766940 1021560 1 0 $X=766940 $Y=1016140
X163 1867 2 1 1827 BUF1 $T=770040 981240 0 180 $X=767560 $Y=975820
X164 155 2 1 1915 BUF1 $T=768180 920760 1 0 $X=768180 $Y=915340
X165 1857 2 1 1913 BUF1 $T=768180 1041720 1 0 $X=768180 $Y=1036300
X166 1867 2 1 1893 BUF1 $T=771280 981240 1 0 $X=771280 $Y=975820
X167 1894 2 1 1871 BUF1 $T=776240 961080 0 180 $X=773760 $Y=955660
X168 1840 2 1 1923 BUF1 $T=778720 1051800 0 180 $X=776240 $Y=1046380
X169 1864 2 1 1894 BUF1 $T=783060 930840 0 180 $X=780580 $Y=925420
X170 1840 2 1 1925 BUF1 $T=780580 1031640 0 0 $X=780580 $Y=1031260
X171 1894 2 1 1950 BUF1 $T=783060 951000 0 0 $X=783060 $Y=950620
X172 1940 2 1 1933 BUF1 $T=784300 951000 1 0 $X=784300 $Y=945580
X173 1913 2 1 1944 BUF1 $T=786780 1051800 1 0 $X=786780 $Y=1046380
X174 1864 2 1 1968 BUF1 $T=791740 920760 0 0 $X=791740 $Y=920380
X175 1913 2 1 1865 BUF1 $T=794220 1051800 0 180 $X=791740 $Y=1046380
X176 1966 2 1 1985 BUF1 $T=795460 1051800 0 0 $X=795460 $Y=1051420
X177 1989 2 1 1980 BUF1 $T=797320 991320 0 0 $X=797320 $Y=990940
X178 1913 2 1 2035 BUF1 $T=798560 1051800 1 0 $X=798560 $Y=1046380
X179 2034 2 1 1989 BUF1 $T=806620 971160 0 180 $X=804140 $Y=965740
X180 1968 2 1 2034 BUF1 $T=805380 940920 0 0 $X=805380 $Y=940540
X181 2035 2 1 2037 BUF1 $T=806000 1031640 0 0 $X=806000 $Y=1031260
X182 2003 2 1 2078 BUF1 $T=809100 971160 0 0 $X=809100 $Y=970780
X183 2034 2 1 2082 BUF1 $T=810960 951000 0 0 $X=810960 $Y=950620
X184 2034 2 1 2088 BUF1 $T=811580 971160 1 0 $X=811580 $Y=965740
X185 2035 2 1 2054 BUF1 $T=812200 1021560 1 0 $X=812200 $Y=1016140
X186 195 2 1 2110 BUF1 $T=817780 910680 0 0 $X=817780 $Y=910300
X187 2121 2 1 2051 BUF1 $T=834520 940920 0 180 $X=832040 $Y=935500
X188 2110 2 1 2121 BUF1 $T=841960 940920 1 0 $X=841960 $Y=935500
X189 216 2 1 209 BUF1 $T=845060 910680 0 180 $X=842580 $Y=905260
X190 2110 2 1 2129 BUF1 $T=842580 930840 1 0 $X=842580 $Y=925420
X191 222 2 1 2136 BUF1 $T=850020 900600 0 0 $X=850020 $Y=900220
X192 2154 2 1 2139 BUF1 $T=859320 920760 1 180 $X=856840 $Y=920380
X193 2134 2 1 2158 BUF1 $T=859320 920760 0 0 $X=859320 $Y=920380
X194 2144 2 1 2163 BUF1 $T=866760 910680 0 0 $X=866760 $Y=910300
X195 2154 2 1 2174 BUF1 $T=870480 940920 1 0 $X=870480 $Y=935500
X196 2149 2 1 2194 BUF1 $T=884740 930840 0 0 $X=884740 $Y=930460
X197 8 6 5 2 1 294 QDFFRBN $T=366420 900600 1 180 $X=354640 $Y=900220
X198 304 6 5 2 1 295 QDFFRBN $T=367660 910680 1 180 $X=355880 $Y=910300
X199 306 6 5 2 1 296 QDFFRBN $T=368280 920760 1 180 $X=356500 $Y=920380
X200 298 6 303 2 1 313 QDFFRBN $T=362080 930840 0 0 $X=362080 $Y=930460
X201 312 6 303 2 1 297 QDFFRBN $T=373860 951000 1 180 $X=362080 $Y=950620
X202 299 6 303 2 1 314 QDFFRBN $T=362700 940920 0 0 $X=362700 $Y=940540
X203 309 6 323 2 1 331 QDFFRBN $T=370140 910680 0 0 $X=370140 $Y=910300
X204 10 6 323 2 1 15 QDFFRBN $T=370760 900600 0 0 $X=370760 $Y=900220
X205 328 6 5 2 1 310 QDFFRBN $T=382540 920760 1 180 $X=370760 $Y=920380
X206 315 6 324 2 1 334 QDFFRBN $T=371380 971160 0 0 $X=371380 $Y=970780
X207 316 6 303 2 1 339 QDFFRBN $T=372620 940920 1 0 $X=372620 $Y=935500
X208 317 6 303 2 1 337 QDFFRBN $T=372620 951000 1 0 $X=372620 $Y=945580
X209 319 6 324 2 1 338 QDFFRBN $T=372620 961080 0 0 $X=372620 $Y=960700
X210 321 6 335 2 1 348 QDFFRBN $T=375720 981240 1 0 $X=375720 $Y=975820
X211 352 340 343 2 1 332 QDFFRBN $T=394320 991320 1 180 $X=382540 $Y=990940
X212 344 6 335 2 1 379 QDFFRBN $T=385640 951000 0 0 $X=385640 $Y=950620
X213 345 6 356 2 1 382 QDFFRBN $T=386260 961080 0 0 $X=386260 $Y=960700
X214 346 6 372 2 1 380 QDFFRBN $T=386260 971160 0 0 $X=386260 $Y=970780
X215 347 6 372 2 1 381 QDFFRBN $T=386260 981240 0 0 $X=386260 $Y=980860
X216 351 6 323 2 1 375 QDFFRBN $T=387500 910680 0 0 $X=387500 $Y=910300
X217 357 6 378 2 1 354 QDFFRBN $T=389360 920760 0 0 $X=389360 $Y=920380
X218 355 6 378 2 1 391 QDFFRBN $T=389360 930840 1 0 $X=389360 $Y=925420
X219 359 6 378 2 1 383 QDFFRBN $T=389980 940920 1 0 $X=389980 $Y=935500
X220 342 6 323 2 1 395 QDFFRBN $T=390600 900600 0 0 $X=390600 $Y=900220
X221 368 340 343 2 1 408 QDFFRBN $T=394940 991320 0 0 $X=394940 $Y=990940
X222 384 6 372 2 1 411 QDFFRBN $T=399280 971160 0 0 $X=399280 $Y=970780
X223 387 6 356 2 1 416 QDFFRBN $T=399900 951000 1 0 $X=399900 $Y=945580
X224 402 6 356 2 1 385 QDFFRBN $T=411680 961080 0 180 $X=399900 $Y=955660
X225 422 6 21 2 1 389 QDFFRBN $T=413540 910680 0 180 $X=401760 $Y=905260
X226 420 6 378 2 1 392 QDFFRBN $T=413540 920760 0 180 $X=401760 $Y=915340
X227 423 6 378 2 1 393 QDFFRBN $T=413540 920760 1 180 $X=401760 $Y=920380
X228 396 340 407 2 1 427 QDFFRBN $T=401760 1031640 0 0 $X=401760 $Y=1031260
X229 410 6 378 2 1 397 QDFFRBN $T=414160 940920 0 180 $X=402380 $Y=935500
X230 415 340 407 2 1 390 QDFFRBN $T=414160 1021560 0 180 $X=402380 $Y=1016140
X231 399 340 407 2 1 433 QDFFRBN $T=403000 1031640 1 0 $X=403000 $Y=1026220
X232 400 6 21 2 1 437 QDFFRBN $T=404240 900600 0 0 $X=404240 $Y=900220
X233 431 6 361 2 1 405 QDFFRBN $T=418500 1001400 0 180 $X=406720 $Y=995980
X234 412 340 361 2 1 450 QDFFRBN $T=407960 1011480 1 0 $X=407960 $Y=1006060
X235 429 6 356 2 1 463 QDFFRBN $T=413540 951000 1 0 $X=413540 $Y=945580
X236 441 340 407 2 1 479 QDFFRBN $T=416020 1021560 1 0 $X=416020 $Y=1016140
X237 447 6 470 2 1 459 QDFFRBN $T=417260 930840 1 0 $X=417260 $Y=925420
X238 448 6 460 2 1 472 QDFFRBN $T=417880 991320 1 0 $X=417880 $Y=985900
X239 430 6 460 2 1 480 QDFFRBN $T=418500 971160 0 0 $X=418500 $Y=970780
X240 434 6 453 2 1 492 QDFFRBN $T=419120 961080 1 0 $X=419120 $Y=955660
X241 455 6 470 2 1 486 QDFFRBN $T=419740 920760 1 0 $X=419740 $Y=915340
X242 456 340 401 2 1 496 QDFFRBN $T=419740 1031640 0 0 $X=419740 $Y=1031260
X243 474 340 361 2 1 457 QDFFRBN $T=432760 1011480 0 180 $X=420980 $Y=1006060
X244 442 340 401 2 1 464 QDFFRBN $T=420980 1041720 1 0 $X=420980 $Y=1036300
X245 508 28 470 2 1 467 QDFFRBN $T=436480 910680 0 180 $X=424700 $Y=905260
X246 478 28 453 2 1 516 QDFFRBN $T=426560 951000 1 0 $X=426560 $Y=945580
X247 469 340 460 2 1 526 QDFFRBN $T=429040 1001400 1 0 $X=429040 $Y=995980
X248 487 340 510 2 1 522 QDFFRBN $T=429040 1021560 1 0 $X=429040 $Y=1016140
X249 527 28 470 2 1 489 QDFFRBN $T=442060 930840 0 180 $X=430280 $Y=925420
X250 498 340 460 2 1 491 QDFFRBN $T=430900 991320 0 0 $X=430900 $Y=990940
X251 471 340 520 2 1 539 QDFFRBN $T=430900 1051800 1 0 $X=430900 $Y=1046380
X252 502 28 525 2 1 517 QDFFRBN $T=432140 961080 0 0 $X=432140 $Y=960700
X253 504 340 401 2 1 545 QDFFRBN $T=432760 1031640 0 0 $X=432760 $Y=1031260
X254 537 28 470 2 1 501 QDFFRBN $T=445160 920760 0 180 $X=433380 $Y=915340
X255 533 340 510 2 1 579 QDFFRBN $T=442060 1021560 1 0 $X=442060 $Y=1016140
X256 538 28 563 2 1 561 QDFFRBN $T=442680 961080 1 0 $X=442680 $Y=955660
X257 562 340 523 2 1 541 QDFFRBN $T=455080 1011480 0 180 $X=443300 $Y=1006060
X258 547 340 510 2 1 589 QDFFRBN $T=445160 1021560 0 0 $X=445160 $Y=1021180
X259 552 340 576 2 1 590 QDFFRBN $T=445780 1031640 0 0 $X=445780 $Y=1031260
X260 556 28 525 2 1 594 QDFFRBN $T=447020 951000 1 0 $X=447020 $Y=945580
X261 557 28 585 2 1 595 QDFFRBN $T=447020 971160 1 0 $X=447020 $Y=965740
X262 558 340 576 2 1 586 QDFFRBN $T=447640 1041720 0 0 $X=447640 $Y=1041340
X263 566 28 525 2 1 600 QDFFRBN $T=450120 940920 0 0 $X=450120 $Y=940540
X264 570 28 597 2 1 614 QDFFRBN $T=450740 930840 1 0 $X=450740 $Y=925420
X265 571 340 523 2 1 615 QDFFRBN $T=450740 1001400 0 0 $X=450740 $Y=1001020
X266 542 28 597 2 1 568 QDFFRBN $T=451360 910680 0 0 $X=451360 $Y=910300
X267 574 28 597 2 1 616 QDFFRBN $T=451360 920760 1 0 $X=451360 $Y=915340
X268 575 340 601 2 1 617 QDFFRBN $T=451360 1061880 1 0 $X=451360 $Y=1056460
X269 581 340 576 2 1 625 QDFFRBN $T=453840 1041720 1 0 $X=453840 $Y=1036300
X270 636 340 510 2 1 593 QDFFRBN $T=469340 1021560 1 180 $X=457560 $Y=1021180
X271 607 28 622 2 1 630 QDFFRBN $T=460040 951000 1 0 $X=460040 $Y=945580
X272 608 28 585 2 1 654 QDFFRBN $T=460040 971160 1 0 $X=460040 $Y=965740
X273 604 340 523 2 1 652 QDFFRBN $T=460040 1011480 0 0 $X=460040 $Y=1011100
X274 629 340 601 2 1 599 QDFFRBN $T=471820 1061880 1 180 $X=460040 $Y=1061500
X275 653 28 622 2 1 611 QDFFRBN $T=472440 940920 0 180 $X=460660 $Y=935500
X276 587 28 585 2 1 633 QDFFRBN $T=461280 981240 1 0 $X=461280 $Y=975820
X277 612 340 585 2 1 639 QDFFRBN $T=461280 991320 1 0 $X=461280 $Y=985900
X278 635 340 523 2 1 619 QDFFRBN $T=474920 1001400 1 180 $X=463140 $Y=1001020
X279 640 28 597 2 1 621 QDFFRBN $T=475540 930840 0 180 $X=463760 $Y=925420
X280 618 28 37 2 1 655 QDFFRBN $T=466860 900600 0 0 $X=466860 $Y=900220
X281 631 28 597 2 1 674 QDFFRBN $T=466860 920760 1 0 $X=466860 $Y=915340
X282 632 28 672 2 1 676 QDFFRBN $T=466860 961080 1 0 $X=466860 $Y=955660
X283 642 340 585 2 1 689 QDFFRBN $T=468100 991320 0 0 $X=468100 $Y=990940
X284 637 340 696 2 1 646 QDFFRBN $T=472440 1021560 0 0 $X=472440 $Y=1021180
X285 716 28 661 2 1 663 QDFFRBN $T=485460 920760 1 180 $X=473680 $Y=920380
X286 666 28 622 2 1 707 QDFFRBN $T=473680 940920 1 0 $X=473680 $Y=935500
X287 667 340 696 2 1 708 QDFFRBN $T=473680 1031640 1 0 $X=473680 $Y=1026220
X288 644 340 601 2 1 711 QDFFRBN $T=474300 1051800 0 0 $X=474300 $Y=1051420
X289 671 340 601 2 1 700 QDFFRBN $T=474300 1061880 0 0 $X=474300 $Y=1061500
X290 678 28 702 2 1 705 QDFFRBN $T=475540 981240 1 0 $X=475540 $Y=975820
X291 680 28 661 2 1 723 QDFFRBN $T=476160 910680 0 0 $X=476160 $Y=910300
X292 683 28 661 2 1 729 QDFFRBN $T=477400 930840 0 0 $X=477400 $Y=930460
X293 681 28 702 2 1 728 QDFFRBN $T=477400 971160 0 0 $X=477400 $Y=970780
X294 685 28 672 2 1 730 QDFFRBN $T=478020 951000 0 0 $X=478020 $Y=950620
X295 688 28 702 2 1 736 QDFFRBN $T=478640 961080 0 0 $X=478640 $Y=960700
X296 697 340 733 2 1 742 QDFFRBN $T=481120 991320 0 0 $X=481120 $Y=990940
X297 698 340 601 2 1 740 QDFFRBN $T=482360 1061880 1 0 $X=482360 $Y=1056460
X298 752 28 704 2 1 713 QDFFRBN $T=497240 910680 0 180 $X=485460 $Y=905260
X299 717 28 622 2 1 765 QDFFRBN $T=485460 940920 0 0 $X=485460 $Y=940540
X300 722 340 746 2 1 773 QDFFRBN $T=487320 1031640 1 0 $X=487320 $Y=1026220
X301 731 340 733 2 1 780 QDFFRBN $T=488560 991320 1 0 $X=488560 $Y=985900
X302 734 28 702 2 1 771 QDFFRBN $T=489180 981240 1 0 $X=489180 $Y=975820
X303 741 46 702 2 1 781 QDFFRBN $T=491660 961080 1 0 $X=491660 $Y=955660
X304 743 46 702 2 1 784 QDFFRBN $T=492280 951000 0 0 $X=492280 $Y=950620
X305 751 340 733 2 1 786 QDFFRBN $T=493520 1001400 1 0 $X=493520 $Y=995980
X306 776 49 47 2 1 754 QDFFRBN $T=506540 910680 1 180 $X=494760 $Y=910300
X307 725 340 750 2 1 798 QDFFRBN $T=494760 1051800 1 0 $X=494760 $Y=1046380
X308 761 46 47 2 1 791 QDFFRBN $T=496000 930840 0 0 $X=496000 $Y=930460
X309 755 340 792 2 1 794 QDFFRBN $T=496000 981240 0 0 $X=496000 $Y=980860
X310 800 46 746 2 1 764 QDFFRBN $T=508400 1011480 1 180 $X=496620 $Y=1011100
X311 766 340 42 2 1 808 QDFFRBN $T=496620 1071960 0 0 $X=496620 $Y=1071580
X312 770 46 750 2 1 821 QDFFRBN $T=497240 1041720 1 0 $X=497240 $Y=1036300
X313 775 46 47 2 1 824 QDFFRBN $T=499100 940920 1 0 $X=499100 $Y=935500
X314 785 340 733 2 1 827 QDFFRBN $T=502820 991320 1 0 $X=502820 $Y=985900
X315 828 49 47 2 1 788 QDFFRBN $T=515220 910680 0 180 $X=503440 $Y=905260
X316 817 49 792 2 1 796 QDFFRBN $T=517080 940920 1 180 $X=505300 $Y=940540
X317 790 46 792 2 1 831 QDFFRBN $T=505300 951000 1 0 $X=505300 $Y=945580
X318 777 340 792 2 1 834 QDFFRBN $T=505300 981240 1 0 $X=505300 $Y=975820
X319 806 46 42 2 1 846 QDFFRBN $T=507160 1061880 0 0 $X=507160 $Y=1061500
X320 809 49 856 2 1 869 QDFFRBN $T=512120 920760 1 0 $X=512120 $Y=915340
X321 833 46 792 2 1 879 QDFFRBN $T=514600 961080 1 0 $X=514600 $Y=955660
X322 829 46 871 2 1 882 QDFFRBN $T=515840 971160 0 0 $X=515840 $Y=970780
X323 839 49 874 2 1 884 QDFFRBN $T=516460 930840 0 0 $X=516460 $Y=930460
X324 842 49 874 2 1 887 QDFFRBN $T=517080 940920 0 0 $X=517080 $Y=940540
X325 849 49 856 2 1 897 QDFFRBN $T=518320 910680 1 0 $X=518320 $Y=905260
X326 812 49 856 2 1 845 QDFFRBN $T=518940 920760 0 0 $X=518940 $Y=920380
X327 852 46 871 2 1 890 QDFFRBN $T=518940 981240 1 0 $X=518940 $Y=975820
X328 853 46 871 2 1 893 QDFFRBN $T=518940 991320 1 0 $X=518940 $Y=985900
X329 855 46 843 2 1 880 QDFFRBN $T=520800 1021560 1 0 $X=520800 $Y=1016140
X330 876 46 891 2 1 927 QDFFRBN $T=524520 1061880 0 0 $X=524520 $Y=1061500
X331 875 46 792 2 1 929 QDFFRBN $T=527000 961080 0 0 $X=527000 $Y=960700
X332 883 46 894 2 1 928 QDFFRBN $T=527000 1011480 1 0 $X=527000 $Y=1006060
X333 896 46 843 2 1 934 QDFFRBN $T=530100 1031640 0 0 $X=530100 $Y=1031260
X334 898 49 931 2 1 942 QDFFRBN $T=530720 940920 0 0 $X=530720 $Y=940540
X335 903 49 917 2 1 945 QDFFRBN $T=531960 910680 1 0 $X=531960 $Y=905260
X336 907 46 940 2 1 957 QDFFRBN $T=533820 981240 1 0 $X=533820 $Y=975820
X337 889 46 894 2 1 948 QDFFRBN $T=533820 1021560 1 0 $X=533820 $Y=1016140
X338 919 46 891 2 1 962 QDFFRBN $T=535060 1061880 1 0 $X=535060 $Y=1056460
X339 918 49 917 2 1 958 QDFFRBN $T=535680 920760 1 0 $X=535680 $Y=915340
X340 923 46 955 2 1 959 QDFFRBN $T=536300 1031640 1 0 $X=536300 $Y=1026220
X341 61 49 917 2 1 62 QDFFRBN $T=536920 900600 0 0 $X=536920 $Y=900220
X342 922 46 940 2 1 970 QDFFRBN $T=537540 971160 0 0 $X=537540 $Y=970780
X343 935 46 967 2 1 976 QDFFRBN $T=539400 940920 1 0 $X=539400 $Y=935500
X344 938 46 955 2 1 984 QDFFRBN $T=540020 1041720 1 0 $X=540020 $Y=1036300
X345 937 46 894 2 1 985 QDFFRBN $T=540640 1011480 1 0 $X=540640 $Y=1006060
X346 944 46 894 2 1 991 QDFFRBN $T=541880 1011480 0 0 $X=541880 $Y=1011100
X347 951 46 940 2 1 979 QDFFRBN $T=543120 991320 1 0 $X=543120 $Y=985900
X348 956 49 917 2 1 1001 QDFFRBN $T=544980 910680 1 0 $X=544980 $Y=905260
X349 963 46 967 2 1 1010 QDFFRBN $T=546220 940920 0 0 $X=546220 $Y=940540
X350 973 46 955 2 1 1023 QDFFRBN $T=549320 1031640 1 0 $X=549320 $Y=1026220
X351 974 46 955 2 1 1024 QDFFRBN $T=549320 1031640 0 0 $X=549320 $Y=1031260
X352 964 46 1013 2 1 996 QDFFRBN $T=549320 1051800 0 0 $X=549320 $Y=1051420
X353 975 46 1013 2 1 1018 QDFFRBN $T=549320 1061880 1 0 $X=549320 $Y=1056460
X354 986 49 931 2 1 1030 QDFFRBN $T=551800 920760 1 0 $X=551800 $Y=915340
X355 990 46 940 2 1 1014 QDFFRBN $T=552420 981240 0 0 $X=552420 $Y=980860
X356 1036 46 1012 2 1 994 QDFFRBN $T=566060 1011480 1 180 $X=554280 $Y=1011100
X357 1006 46 939 2 1 1040 QDFFRBN $T=556140 951000 0 0 $X=556140 $Y=950620
X358 1015 49 64 2 1 1062 QDFFRBN $T=558000 910680 1 0 $X=558000 $Y=905260
X359 1016 49 1045 2 1 1063 QDFFRBN $T=558000 910680 0 0 $X=558000 $Y=910300
X360 1017 46 1027 2 1 1057 QDFFRBN $T=558000 971160 1 0 $X=558000 $Y=965740
X361 1021 1026 967 2 1 1068 QDFFRBN $T=559240 940920 0 0 $X=559240 $Y=940540
X362 1033 46 1069 2 1 1056 QDFFRBN $T=562340 1061880 1 0 $X=562340 $Y=1056460
X363 1037 46 1013 2 1 1086 QDFFRBN $T=562960 1031640 0 0 $X=562960 $Y=1031260
X364 1039 49 1076 2 1 1088 QDFFRBN $T=563580 930840 0 0 $X=563580 $Y=930460
X365 1044 63 1084 2 1 1097 QDFFRBN $T=565440 991320 1 0 $X=565440 $Y=985900
X366 1072 63 1012 2 1 1047 QDFFRBN $T=577840 1001400 1 180 $X=566060 $Y=1001020
X367 1054 46 1012 2 1 1107 QDFFRBN $T=566680 1011480 0 0 $X=566680 $Y=1011100
X368 1104 1026 1061 2 1 1055 QDFFRBN $T=579700 961080 0 180 $X=567920 $Y=955660
X369 1059 46 367 2 1 1111 QDFFRBN $T=567920 1051800 0 0 $X=567920 $Y=1051420
X370 1105 1026 1061 2 1 1064 QDFFRBN $T=580940 961080 1 180 $X=569160 $Y=960700
X371 1074 49 1045 2 1 1124 QDFFRBN $T=571020 910680 1 0 $X=571020 $Y=905260
X372 1075 49 1045 2 1 1125 QDFFRBN $T=571020 910680 0 0 $X=571020 $Y=910300
X373 1079 1026 1117 2 1 1116 QDFFRBN $T=572880 940920 0 0 $X=572880 $Y=940540
X374 1119 63 1084 2 1 1090 QDFFRBN $T=586520 1001400 0 180 $X=574740 $Y=995980
X375 1099 1026 1076 2 1 1141 QDFFRBN $T=576600 940920 1 0 $X=576600 $Y=935500
X376 1095 63 1084 2 1 1131 QDFFRBN $T=576600 1011480 1 0 $X=576600 $Y=1006060
X377 1091 63 1069 2 1 1143 QDFFRBN $T=576600 1041720 0 0 $X=576600 $Y=1041340
X378 1087 63 1142 2 1 1133 QDFFRBN $T=579700 1021560 0 0 $X=579700 $Y=1021180
X379 1115 63 1142 2 1 1155 QDFFRBN $T=579700 1031640 1 0 $X=579700 $Y=1026220
X380 1098 1026 1076 2 1 1161 QDFFRBN $T=580940 930840 0 0 $X=580940 $Y=930460
X381 1120 63 1069 2 1 1137 QDFFRBN $T=580940 1051800 1 0 $X=580940 $Y=1046380
X382 1127 63 1149 2 1 1166 QDFFRBN $T=582800 981240 1 0 $X=582800 $Y=975820
X383 1130 49 1045 2 1 1173 QDFFRBN $T=584040 910680 1 0 $X=584040 $Y=905260
X384 1136 63 1069 2 1 1171 QDFFRBN $T=585900 1061880 0 0 $X=585900 $Y=1061500
X385 1138 63 1142 2 1 1186 QDFFRBN $T=586520 1021560 1 0 $X=586520 $Y=1016140
X386 1135 1026 1172 2 1 1189 QDFFRBN $T=587140 961080 1 0 $X=587140 $Y=955660
X387 1140 63 1149 2 1 1190 QDFFRBN $T=587140 1001400 1 0 $X=587140 $Y=995980
X388 1144 1026 1172 2 1 1196 QDFFRBN $T=587760 951000 1 0 $X=587760 $Y=945580
X389 1191 63 1149 2 1 1145 QDFFRBN $T=600160 981240 1 180 $X=588380 $Y=980860
X390 1150 63 1187 2 1 1199 QDFFRBN $T=589620 1041720 0 0 $X=589620 $Y=1041340
X391 1153 63 1187 2 1 1202 QDFFRBN $T=590240 1041720 1 0 $X=590240 $Y=1036300
X392 1179 63 1142 2 1 1158 QDFFRBN $T=603260 1031640 0 180 $X=591480 $Y=1026220
X393 1164 1026 1207 2 1 1221 QDFFRBN $T=594580 920760 0 0 $X=594580 $Y=920380
X394 1180 63 1213 2 1 1228 QDFFRBN $T=595820 1071960 1 0 $X=595820 $Y=1066540
X395 1245 63 1069 2 1 1183 QDFFRBN $T=608220 1061880 0 180 $X=596440 $Y=1056460
X396 1165 1026 1217 2 1 1233 QDFFRBN $T=597060 971160 1 0 $X=597060 $Y=965740
X397 1185 63 1149 2 1 1236 QDFFRBN $T=597060 1011480 1 0 $X=597060 $Y=1006060
X398 1203 1026 1172 2 1 1194 QDFFRBN $T=611320 961080 0 180 $X=599540 $Y=955660
X399 1197 63 1235 2 1 1248 QDFFRBN $T=600160 1021560 0 0 $X=600160 $Y=1021180
X400 1206 63 1235 2 1 1251 QDFFRBN $T=602020 1031640 0 0 $X=602020 $Y=1031260
X401 1220 1026 1172 2 1 1262 QDFFRBN $T=605120 951000 1 0 $X=605120 $Y=945580
X402 1258 63 1237 2 1 1219 QDFFRBN $T=617520 1001400 1 180 $X=605740 $Y=1001020
X403 1204 63 1235 2 1 1268 QDFFRBN $T=606360 1021560 1 0 $X=606360 $Y=1016140
X404 1229 1026 1207 2 1 1256 QDFFRBN $T=606980 940920 1 0 $X=606980 $Y=935500
X405 1230 63 1237 2 1 1274 QDFFRBN $T=606980 991320 0 0 $X=606980 $Y=990940
X406 1205 74 1259 2 1 86 QDFFRBN $T=607600 900600 0 0 $X=607600 $Y=900220
X407 1231 74 1259 2 1 1272 QDFFRBN $T=607600 920760 1 0 $X=607600 $Y=915340
X408 1240 1026 1217 2 1 1271 QDFFRBN $T=608840 961080 0 0 $X=608840 $Y=960700
X409 85 63 1213 2 1 80 QDFFRBN $T=620620 1071960 1 180 $X=608840 $Y=1071580
X410 1226 63 1187 2 1 1286 QDFFRBN $T=610700 1051800 1 0 $X=610700 $Y=1046380
X411 1246 63 1213 2 1 1292 QDFFRBN $T=611320 1061880 1 0 $X=611320 $Y=1056460
X412 1275 63 1235 2 1 1253 QDFFRBN $T=625580 1031640 1 180 $X=613800 $Y=1031260
X413 1257 63 1237 2 1 1310 QDFFRBN $T=615040 1001400 1 0 $X=615040 $Y=995980
X414 1261 63 1235 2 1 1306 QDFFRBN $T=615660 1021560 0 0 $X=615660 $Y=1021180
X415 1263 63 1296 2 1 1312 QDFFRBN $T=616280 991320 1 0 $X=616280 $Y=985900
X416 1269 63 1213 2 1 1317 QDFFRBN $T=617520 1061880 0 0 $X=617520 $Y=1061500
X417 1270 1026 1305 2 1 1308 QDFFRBN $T=618140 951000 1 0 $X=618140 $Y=945580
X418 1304 63 1237 2 1 1273 QDFFRBN $T=630540 1001400 1 180 $X=618760 $Y=1001020
X419 1282 74 1259 2 1 93 QDFFRBN $T=620620 900600 0 0 $X=620620 $Y=900220
X420 1283 1026 1305 2 1 1319 QDFFRBN $T=620620 940920 1 0 $X=620620 $Y=935500
X421 1284 1026 1217 2 1 1313 QDFFRBN $T=620620 981240 1 0 $X=620620 $Y=975820
X422 87 63 1213 2 1 92 QDFFRBN $T=621240 1071960 0 0 $X=621240 $Y=1071580
X423 1316 63 1187 2 1 1290 QDFFRBN $T=634260 1051800 0 180 $X=622480 $Y=1046380
X424 1329 74 1259 2 1 1285 QDFFRBN $T=634880 910680 1 180 $X=623100 $Y=910300
X425 1287 74 1259 2 1 1341 QDFFRBN $T=623720 920760 1 0 $X=623720 $Y=915340
X426 1327 63 1235 2 1 1302 QDFFRBN $T=637360 1031640 1 180 $X=625580 $Y=1031260
X427 89 74 1300 2 1 1359 QDFFRBN $T=628680 910680 1 0 $X=628680 $Y=905260
X428 1297 1026 1345 2 1 1356 QDFFRBN $T=628680 930840 1 0 $X=628680 $Y=925420
X429 1318 1026 1345 2 1 1348 QDFFRBN $T=628680 940920 0 0 $X=628680 $Y=940540
X430 1320 1026 1350 2 1 1342 QDFFRBN $T=629300 981240 0 0 $X=629300 $Y=980860
X431 1323 63 1350 2 1 1368 QDFFRBN $T=631160 1001400 0 0 $X=631160 $Y=1001020
X432 1375 63 1340 2 1 1326 QDFFRBN $T=644180 1061880 0 180 $X=632400 $Y=1056460
X433 1330 1026 1350 2 1 1367 QDFFRBN $T=633020 991320 0 0 $X=633020 $Y=990940
X434 1374 1026 1321 2 1 1331 QDFFRBN $T=645420 961080 1 180 $X=633640 $Y=960700
X435 1376 63 91 2 1 1333 QDFFRBN $T=645420 1071960 1 180 $X=633640 $Y=1071580
X436 1336 63 1340 2 1 1382 QDFFRBN $T=634260 1051800 1 0 $X=634260 $Y=1046380
X437 1349 1026 1350 2 1 1396 QDFFRBN $T=636740 981240 1 0 $X=636740 $Y=975820
X438 1352 63 1384 2 1 1365 QDFFRBN $T=637360 1031640 0 0 $X=637360 $Y=1031260
X439 1354 1026 1345 2 1 1392 QDFFRBN $T=637980 930840 0 0 $X=637980 $Y=930460
X440 1378 74 1345 2 1 1362 QDFFRBN $T=652240 920760 1 180 $X=640460 $Y=920380
X441 99 74 94 2 1 103 QDFFRBN $T=642940 900600 0 0 $X=642940 $Y=900220
X442 1364 74 94 2 1 1418 QDFFRBN $T=642940 910680 1 0 $X=642940 $Y=905260
X443 1373 1026 1345 2 1 1419 QDFFRBN $T=642940 940920 0 0 $X=642940 $Y=940540
X444 1399 1026 1350 2 1 1370 QDFFRBN $T=654720 991320 0 180 $X=642940 $Y=985900
X445 1405 63 1350 2 1 1371 QDFFRBN $T=654720 1001400 1 180 $X=642940 $Y=1001020
X446 1389 74 94 2 1 1433 QDFFRBN $T=646040 910680 0 0 $X=646040 $Y=910300
X447 1429 63 1340 2 1 1388 QDFFRBN $T=657820 1061880 0 180 $X=646040 $Y=1056460
X448 1390 63 91 2 1 1435 QDFFRBN $T=646040 1071960 0 0 $X=646040 $Y=1071580
X449 1432 102 1384 2 1 1391 QDFFRBN $T=658440 1051800 0 180 $X=646660 $Y=1046380
X450 1393 102 1434 2 1 1445 QDFFRBN $T=649140 1021560 1 0 $X=649140 $Y=1016140
X451 1431 102 1384 2 1 1401 QDFFRBN $T=660920 1031640 1 180 $X=649140 $Y=1031260
X452 1407 1026 1321 2 1 1436 QDFFRBN $T=650380 951000 0 0 $X=650380 $Y=950620
X453 1422 74 1438 2 1 1461 QDFFRBN $T=654720 930840 1 0 $X=654720 $Y=925420
X454 1423 63 1454 2 1 1468 QDFFRBN $T=654720 1001400 0 0 $X=654720 $Y=1001020
X455 1416 63 1454 2 1 1421 QDFFRBN $T=655340 991320 0 0 $X=655340 $Y=990940
X456 1427 63 1417 2 1 1472 QDFFRBN $T=655340 1061880 0 0 $X=655340 $Y=1061500
X457 1442 74 1438 2 1 1476 QDFFRBN $T=658440 920760 1 0 $X=658440 $Y=915340
X458 1447 74 111 2 1 113 QDFFRBN $T=660920 900600 0 0 $X=660920 $Y=900220
X459 1449 102 1434 2 1 1491 QDFFRBN $T=660920 1021560 0 0 $X=660920 $Y=1021180
X460 1485 102 1463 2 1 1446 QDFFRBN $T=672700 1031640 1 180 $X=660920 $Y=1031260
X461 1451 102 1434 2 1 1494 QDFFRBN $T=661540 1011480 0 0 $X=661540 $Y=1011100
X462 1459 1026 1489 2 1 1495 QDFFRBN $T=663400 951000 0 0 $X=663400 $Y=950620
X463 1466 102 1463 2 1 1506 QDFFRBN $T=664020 1041720 0 0 $X=664020 $Y=1041340
X464 1497 102 1417 2 1 1458 QDFFRBN $T=677660 1061880 0 180 $X=665880 $Y=1056460
X465 1511 102 1454 2 1 1470 QDFFRBN $T=678280 1001400 1 180 $X=666500 $Y=1001020
X466 1496 102 1486 2 1 1469 QDFFRBN $T=679520 991320 0 180 $X=667740 $Y=985900
X467 1480 1026 1507 2 1 1523 QDFFRBN $T=668360 930840 1 0 $X=668360 $Y=925420
X468 1524 74 1438 2 1 1481 QDFFRBN $T=681380 910680 1 180 $X=669600 $Y=910300
X469 1484 102 1486 2 1 1526 QDFFRBN $T=669600 981240 0 0 $X=669600 $Y=980860
X470 1528 102 1417 2 1 1479 QDFFRBN $T=682000 1051800 1 180 $X=670220 $Y=1051420
X471 1493 102 121 2 1 1540 QDFFRBN $T=672080 1071960 1 0 $X=672080 $Y=1066540
X472 1499 102 1463 2 1 1544 QDFFRBN $T=673320 1031640 0 0 $X=673320 $Y=1031260
X473 1500 1026 1507 2 1 1547 QDFFRBN $T=673940 930840 0 0 $X=673940 $Y=930460
X474 1501 1026 1489 2 1 1542 QDFFRBN $T=673940 951000 1 0 $X=673940 $Y=945580
X475 1508 1026 1489 2 1 1541 QDFFRBN $T=675800 961080 0 0 $X=675800 $Y=960700
X476 1552 1026 1489 2 1 1509 QDFFRBN $T=688200 951000 1 180 $X=676420 $Y=950620
X477 1536 102 1513 2 1 1510 QDFFRBN $T=688200 1011480 1 180 $X=676420 $Y=1011100
X478 1516 102 1513 2 1 1564 QDFFRBN $T=677660 1011480 1 0 $X=677660 $Y=1006060
X479 1559 102 1463 2 1 1514 QDFFRBN $T=689440 1041720 0 180 $X=677660 $Y=1036300
X480 1517 102 1463 2 1 1563 QDFFRBN $T=677660 1041720 0 0 $X=677660 $Y=1041340
X481 1525 102 1513 2 1 1576 QDFFRBN $T=679520 1001400 1 0 $X=679520 $Y=995980
X482 1527 102 1486 2 1 1568 QDFFRBN $T=680140 991320 1 0 $X=680140 $Y=985900
X483 1551 127 111 2 1 123 QDFFRBN $T=692540 900600 1 180 $X=680760 $Y=900220
X484 1533 1026 1507 2 1 1565 QDFFRBN $T=681380 920760 0 0 $X=681380 $Y=920380
X485 1582 102 1434 2 1 1531 QDFFRBN $T=693160 1021560 0 180 $X=681380 $Y=1016140
X486 1535 1026 1507 2 1 1570 QDFFRBN $T=682000 930840 1 0 $X=682000 $Y=925420
X487 1566 102 121 2 1 1530 QDFFRBN $T=693780 1061880 1 180 $X=682000 $Y=1061500
X488 1550 1026 1585 2 1 1599 QDFFRBN $T=685720 940920 0 0 $X=685720 $Y=940540
X489 1600 102 1463 2 1 1555 QDFFRBN $T=698740 1031640 1 180 $X=686960 $Y=1031260
X490 131 102 1578 2 1 126 QDFFRBN $T=699360 1071960 1 180 $X=687580 $Y=1071580
X491 1604 1026 1489 2 1 1560 QDFFRBN $T=700600 951000 1 180 $X=688820 $Y=950620
X492 1574 1026 1603 2 1 1622 QDFFRBN $T=690060 920760 1 0 $X=690060 $Y=915340
X493 1611 1026 1581 2 1 1571 QDFFRBN $T=701840 961080 1 180 $X=690060 $Y=960700
X494 1575 1026 1581 2 1 1620 QDFFRBN $T=690060 971160 1 0 $X=690060 $Y=965740
X495 1584 102 1585 2 1 1631 QDFFRBN $T=692540 1001400 1 0 $X=692540 $Y=995980
X496 1629 102 1513 2 1 1586 QDFFRBN $T=705560 991320 0 180 $X=693780 $Y=985900
X497 1590 102 1513 2 1 1640 QDFFRBN $T=694400 1011480 0 0 $X=694400 $Y=1011100
X498 1591 102 1624 2 1 1639 QDFFRBN $T=694400 1021560 1 0 $X=694400 $Y=1016140
X499 1592 102 1625 2 1 1638 QDFFRBN $T=694400 1061880 1 0 $X=694400 $Y=1056460
X500 1594 102 1625 2 1 1642 QDFFRBN $T=695020 1061880 0 0 $X=695020 $Y=1061500
X501 1601 102 1624 2 1 1646 QDFFRBN $T=696880 1041720 1 0 $X=696880 $Y=1036300
X502 1647 1583 1617 2 1 1598 QDFFRBN $T=709900 940920 0 180 $X=698120 $Y=935500
X503 1671 102 1585 2 1 1609 QDFFRBN $T=711760 991320 1 180 $X=699980 $Y=990940
X504 1665 102 1578 2 1 1616 QDFFRBN $T=712380 1071960 1 180 $X=700600 $Y=1071580
X505 1628 1026 1666 2 1 1670 QDFFRBN $T=703080 951000 0 0 $X=703080 $Y=950620
X506 1633 1026 1603 2 1 1687 QDFFRBN $T=703700 920760 1 0 $X=703700 $Y=915340
X507 1658 102 1624 2 1 1644 QDFFRBN $T=718580 1021560 0 180 $X=706800 $Y=1016140
X508 1648 1583 1617 2 1 1700 QDFFRBN $T=708040 940920 0 0 $X=708040 $Y=940540
X509 1699 1026 1666 2 1 1650 QDFFRBN $T=720440 961080 0 180 $X=708660 $Y=955660
X510 1663 102 1624 2 1 1716 QDFFRBN $T=710520 1021560 0 0 $X=710520 $Y=1021180
X511 1656 127 1703 2 1 1660 QDFFRBN $T=711760 910680 0 0 $X=711760 $Y=910300
X512 1678 1583 1685 2 1 1662 QDFFRBN $T=723540 971160 1 180 $X=711760 $Y=970780
X513 1668 102 1625 2 1 1655 QDFFRBN $T=724160 1061880 0 180 $X=712380 $Y=1056460
X514 1718 1583 1685 2 1 1680 QDFFRBN $T=726020 981240 0 180 $X=714240 $Y=975820
X515 1695 102 1691 2 1 1674 QDFFRBN $T=726020 1051800 0 180 $X=714240 $Y=1046380
X516 1722 102 130 2 1 1673 QDFFRBN $T=726020 1071960 0 180 $X=714240 $Y=1066540
X517 1717 1583 1603 2 1 1684 QDFFRBN $T=726640 930840 0 180 $X=714860 $Y=925420
X518 1694 102 1732 2 1 1740 QDFFRBN $T=719820 991320 0 0 $X=719820 $Y=990940
X519 1707 102 1732 2 1 1743 QDFFRBN $T=720440 1001400 0 0 $X=720440 $Y=1001020
X520 1710 1026 1666 2 1 1739 QDFFRBN $T=721060 961080 1 0 $X=721060 $Y=955660
X521 1688 147 1685 2 1 1705 QDFFRBN $T=732840 991320 0 180 $X=721060 $Y=985900
X522 1713 1583 1736 2 1 1745 QDFFRBN $T=721680 940920 0 0 $X=721680 $Y=940540
X523 1715 102 1738 2 1 1749 QDFFRBN $T=721680 1051800 0 0 $X=721680 $Y=1051420
X524 1750 127 1703 2 1 141 QDFFRBN $T=734700 900600 1 180 $X=722920 $Y=900220
X525 1692 1583 1736 2 1 1757 QDFFRBN $T=722920 940920 1 0 $X=722920 $Y=935500
X526 1719 102 1744 2 1 1752 QDFFRBN $T=723540 1021560 1 0 $X=723540 $Y=1016140
X527 1723 102 1738 2 1 1772 QDFFRBN $T=724780 1061880 0 0 $X=724780 $Y=1061500
X528 1728 127 1703 2 1 1768 QDFFRBN $T=725400 910680 0 0 $X=725400 $Y=910300
X529 1766 1583 1617 2 1 1725 QDFFRBN $T=737800 930840 1 180 $X=726020 $Y=930460
X530 1751 1583 1685 2 1 1727 QDFFRBN $T=737800 981240 0 180 $X=726020 $Y=975820
X531 1780 147 1734 2 1 1731 QDFFRBN $T=739660 1051800 0 180 $X=727880 $Y=1046380
X532 1788 1583 1759 2 1 1742 QDFFRBN $T=743380 961080 1 180 $X=731600 $Y=960700
X533 1770 147 1732 2 1 1747 QDFFRBN $T=744000 1001400 1 180 $X=732220 $Y=1001020
X534 1741 1583 1785 2 1 1735 QDFFRBN $T=733460 920760 0 0 $X=733460 $Y=920380
X535 1779 1583 1736 2 1 1753 QDFFRBN $T=745240 940920 1 180 $X=733460 $Y=940540
X536 1755 147 1732 2 1 1802 QDFFRBN $T=733460 1001400 1 0 $X=733460 $Y=995980
X537 1799 147 1734 2 1 1754 QDFFRBN $T=745240 1041720 0 180 $X=733460 $Y=1036300
X538 1797 1583 1759 2 1 1758 QDFFRBN $T=746480 961080 0 180 $X=734700 $Y=955660
X539 1809 1583 1685 2 1 1761 QDFFRBN $T=746480 971160 1 180 $X=734700 $Y=970780
X540 1817 127 157 2 1 1775 QDFFRBN $T=750200 910680 0 180 $X=738420 $Y=905260
X541 1787 1583 1785 2 1 1832 QDFFRBN $T=740900 920760 1 0 $X=740900 $Y=915340
X542 1789 147 1756 2 1 1835 QDFFRBN $T=741520 1061880 1 0 $X=741520 $Y=1056460
X543 1794 1583 1736 2 1 1830 QDFFRBN $T=742760 940920 1 0 $X=742760 $Y=935500
X544 1795 147 1732 2 1 1801 QDFFRBN $T=742760 991320 1 0 $X=742760 $Y=985900
X545 1818 147 1806 2 1 1792 QDFFRBN $T=754540 1011480 0 180 $X=742760 $Y=1006060
X546 1812 147 1756 2 1 1790 QDFFRBN $T=754540 1051800 1 180 $X=742760 $Y=1051420
X547 1839 147 1744 2 1 1800 QDFFRBN $T=756400 1031640 0 180 $X=744620 $Y=1026220
X548 1805 1583 1831 2 1 1843 QDFFRBN $T=745240 940920 0 0 $X=745240 $Y=940540
X549 1807 147 1732 2 1 1853 QDFFRBN $T=745860 1001400 0 0 $X=745860 $Y=1001020
X550 1810 147 1840 2 1 1854 QDFFRBN $T=746480 1051800 1 0 $X=746480 $Y=1046380
X551 1811 147 1827 2 1 1856 QDFFRBN $T=747100 981240 0 0 $X=747100 $Y=980860
X552 1837 1583 1827 2 1 1813 QDFFRBN $T=759500 981240 0 180 $X=747720 $Y=975820
X553 1820 1583 1831 2 1 1862 QDFFRBN $T=748960 961080 1 0 $X=748960 $Y=955660
X554 1829 127 1785 2 1 1866 QDFFRBN $T=750820 910680 1 0 $X=750820 $Y=905260
X555 1875 1583 1785 2 1 1821 QDFFRBN $T=762600 920760 1 180 $X=750820 $Y=920380
X556 1834 1583 1831 2 1 1877 QDFFRBN $T=752060 951000 1 0 $X=752060 $Y=945580
X557 1873 147 1806 2 1 1833 QDFFRBN $T=763840 1011480 1 180 $X=752060 $Y=1011100
X558 1836 147 1806 2 1 1884 QDFFRBN $T=753300 1021560 0 0 $X=753300 $Y=1021180
X559 166 127 160 2 1 170 QDFFRBN $T=753920 900600 0 0 $X=753920 $Y=900220
X560 1838 1583 1867 2 1 1886 QDFFRBN $T=753920 971160 0 0 $X=753920 $Y=970780
X561 1878 147 1756 2 1 1841 QDFFRBN $T=766320 1061880 0 180 $X=754540 $Y=1056460
X562 1905 1583 1831 2 1 1844 QDFFRBN $T=767560 951000 1 180 $X=755780 $Y=950620
X563 1891 147 1806 2 1 1845 QDFFRBN $T=767560 1011480 0 180 $X=755780 $Y=1006060
X564 1892 147 164 2 1 1850 QDFFRBN $T=768180 1071960 0 180 $X=756400 $Y=1066540
X565 1870 1583 1831 2 1 1851 QDFFRBN $T=768800 940920 1 180 $X=757020 $Y=940540
X566 1858 147 1893 2 1 1897 QDFFRBN $T=758880 991320 1 0 $X=758880 $Y=985900
X567 1881 147 1840 2 1 1863 QDFFRBN $T=771900 1051800 0 180 $X=760120 $Y=1046380
X568 1910 127 1785 2 1 1874 QDFFRBN $T=774380 910680 0 180 $X=762600 $Y=905260
X569 1909 147 1840 2 1 1876 QDFFRBN $T=775000 1031640 1 180 $X=763220 $Y=1031260
X570 1926 1583 1785 2 1 1879 QDFFRBN $T=775620 920760 1 180 $X=763840 $Y=920380
X571 1888 147 1925 2 1 1918 QDFFRBN $T=765080 1011480 0 0 $X=765080 $Y=1011100
X572 1929 1583 1867 2 1 1896 QDFFRBN $T=779960 971160 1 180 $X=768180 $Y=970780
X573 1900 147 1923 2 1 1946 QDFFRBN $T=768180 1041720 0 0 $X=768180 $Y=1041340
X574 1902 1583 1933 2 1 1943 QDFFRBN $T=768800 930840 0 0 $X=768800 $Y=930460
X575 1947 147 1923 2 1 1903 QDFFRBN $T=781200 1061880 0 180 $X=769420 $Y=1056460
X576 1948 147 164 2 1 1904 QDFFRBN $T=781200 1071960 0 180 $X=769420 $Y=1066540
X577 1911 1583 1940 2 1 1953 QDFFRBN $T=770660 951000 0 0 $X=770660 $Y=950620
X578 1916 1583 1893 2 1 1958 QDFFRBN $T=771280 981240 0 0 $X=771280 $Y=980860
X579 1921 127 19 2 1 1961 QDFFRBN $T=771900 910680 0 0 $X=771900 $Y=910300
X580 1935 147 1925 2 1 1920 QDFFRBN $T=783680 1031640 0 180 $X=771900 $Y=1026220
X581 1930 1583 1867 2 1 1975 QDFFRBN $T=775620 981240 1 0 $X=775620 $Y=975820
X582 1960 147 1925 2 1 1934 QDFFRBN $T=788640 1011480 1 180 $X=776860 $Y=1011100
X583 1979 1583 1940 2 1 1937 QDFFRBN $T=789260 961080 0 180 $X=777480 $Y=955660
X584 1939 147 1925 2 1 1987 QDFFRBN $T=778100 1021560 0 0 $X=778100 $Y=1021180
X585 1956 1583 1933 2 1 2005 QDFFRBN $T=781820 930840 0 0 $X=781820 $Y=930460
X586 2002 147 1966 2 1 1949 QDFFRBN $T=793600 1041720 1 180 $X=781820 $Y=1041340
X587 1969 147 1966 2 1 2014 QDFFRBN $T=784920 1041720 1 0 $X=784920 $Y=1036300
X588 1997 147 1985 2 1 1967 QDFFRBN $T=797940 1061880 0 180 $X=786160 $Y=1056460
X589 1978 1583 1940 2 1 2029 QDFFRBN $T=787400 951000 1 0 $X=787400 $Y=945580
X590 1981 147 1985 2 1 2027 QDFFRBN $T=787400 1061880 0 0 $X=787400 $Y=1061500
X591 1983 1583 2003 2 1 2010 QDFFRBN $T=788020 971160 0 0 $X=788020 $Y=970780
X592 1986 147 2019 2 1 2018 QDFFRBN $T=789260 1001400 0 0 $X=789260 $Y=1001020
X593 1984 147 2019 2 1 2040 QDFFRBN $T=789260 1011480 0 0 $X=789260 $Y=1011100
X594 1990 1583 1940 2 1 2036 QDFFRBN $T=790500 961080 1 0 $X=790500 $Y=955660
X595 1996 147 2003 2 1 2043 QDFFRBN $T=791120 991320 1 0 $X=791120 $Y=985900
X596 2004 147 2033 2 1 2048 QDFFRBN $T=792360 1031640 1 0 $X=792360 $Y=1026220
X597 2020 1583 2051 2 1 2047 QDFFRBN $T=796700 930840 0 0 $X=796700 $Y=930460
X598 2061 147 2019 2 1 2017 QDFFRBN $T=808480 1011480 0 180 $X=796700 $Y=1006060
X599 2021 1583 2051 2 1 2068 QDFFRBN $T=797320 940920 1 0 $X=797320 $Y=935500
X600 2042 147 1985 2 1 2031 QDFFRBN $T=810960 1061880 0 180 $X=799180 $Y=1056460
X601 2046 1583 2078 2 1 2083 QDFFRBN $T=803520 961080 1 0 $X=803520 $Y=955660
X602 2065 147 2033 2 1 2044 QDFFRBN $T=815920 1041720 1 180 $X=804140 $Y=1041340
X603 2079 147 2019 2 1 2057 QDFFRBN $T=818400 991320 1 180 $X=806620 $Y=990940
X604 2030 127 195 2 1 2059 QDFFRBN $T=819020 910680 0 180 $X=807240 $Y=905260
X605 2056 147 1966 2 1 2105 QDFFRBN $T=808480 1051800 0 0 $X=808480 $Y=1051420
X606 2076 147 2101 2 1 2103 QDFFRBN $T=810960 1011480 1 0 $X=810960 $Y=1006060
X607 2077 147 1966 2 1 2109 QDFFRBN $T=810960 1051800 1 0 $X=810960 $Y=1046380
X608 2075 1583 2110 2 1 199 QDFFRBN $T=814060 920760 0 0 $X=814060 $Y=920380
X609 2063 1583 2051 2 1 2081 QDFFRBN $T=814060 930840 1 0 $X=814060 $Y=925420
X610 2060 1583 2110 2 1 202 QDFFRBN $T=814680 920760 1 0 $X=814680 $Y=915340
X611 2090 1583 2051 2 1 2115 QDFFRBN $T=814680 930840 0 0 $X=814680 $Y=930460
X612 2100 1583 2078 2 1 2085 QDFFRBN $T=827700 971160 1 180 $X=815920 $Y=970780
X613 2112 147 2101 2 1 2095 QDFFRBN $T=827700 1001400 0 180 $X=815920 $Y=995980
X614 2097 147 2033 2 1 2118 QDFFRBN $T=816540 1021560 0 0 $X=816540 $Y=1021180
X615 2080 147 2033 2 1 2119 QDFFRBN $T=816540 1031640 0 0 $X=816540 $Y=1031260
X616 2058 127 200 2 1 206 QDFFRBN $T=820260 910680 1 0 $X=820260 $Y=905260
X617 2094 1583 2078 2 1 2123 QDFFRBN $T=820880 961080 0 0 $X=820880 $Y=960700
X618 2108 147 2101 2 1 2124 QDFFRBN $T=820880 1001400 0 0 $X=820880 $Y=1001020
X619 2084 1583 2121 2 1 2126 QDFFRBN $T=822120 940920 0 0 $X=822120 $Y=940540
X620 2099 1583 2121 2 1 2127 QDFFRBN $T=822120 951000 1 0 $X=822120 $Y=945580
X621 2111 1583 2078 2 1 2102 QDFFRBN $T=822120 961080 1 0 $X=822120 $Y=955660
X622 2113 1583 2078 2 1 2128 QDFFRBN $T=823360 981240 1 0 $X=823360 $Y=975820
X623 201 1583 2129 2 1 213 QDFFRBN $T=826460 910680 0 0 $X=826460 $Y=910300
X624 2116 147 2101 2 1 2130 QDFFRBN $T=826460 1011480 1 0 $X=826460 $Y=1006060
X625 2066 1583 2110 2 1 210 QDFFRBN $T=827080 920760 0 0 $X=827080 $Y=920380
X626 1711 1583 2110 2 1 215 QDFFRBN $T=827700 930840 1 0 $X=827700 $Y=925420
X627 2032 1583 2129 2 1 212 QDFFRBN $T=828320 920760 1 0 $X=828320 $Y=915340
X628 2120 147 2101 2 1 2131 QDFFRBN $T=829560 1001400 1 0 $X=829560 $Y=995980
X629 2049 1583 2121 2 1 2152 QDFFRBN $T=835760 940920 0 0 $X=835760 $Y=940540
X630 2067 1583 2121 2 1 2141 QDFFRBN $T=835760 951000 1 0 $X=835760 $Y=945580
X631 295 2 301 1 INV1S $T=363320 920760 1 0 $X=363320 $Y=915340
X632 294 2 9 1 INV1S $T=367660 900600 0 0 $X=367660 $Y=900220
X633 313 2 302 1 INV1S $T=370760 940920 0 180 $X=369520 $Y=935500
X634 296 2 300 1 INV1S $T=370140 930840 1 0 $X=370140 $Y=925420
X635 314 2 307 1 INV1S $T=371380 951000 0 180 $X=370140 $Y=945580
X636 297 2 311 1 INV1S $T=370140 961080 0 0 $X=370140 $Y=960700
X637 12 2 324 1 INV1S $T=377580 1071960 0 0 $X=377580 $Y=1071580
X638 331 2 325 1 INV1S $T=383160 910680 0 0 $X=383160 $Y=910300
X639 310 2 336 1 INV1S $T=383160 920760 0 0 $X=383160 $Y=920380
X640 338 2 322 1 INV1S $T=384400 961080 0 180 $X=383160 $Y=955660
X641 337 2 327 1 INV1S $T=383780 951000 0 0 $X=383780 $Y=950620
X642 334 2 320 1 INV1S $T=385020 971160 1 0 $X=385020 $Y=965740
X643 12 2 350 1 INV1S $T=385020 1051800 0 0 $X=385020 $Y=1051420
X644 339 2 341 1 INV1S $T=385640 940920 1 0 $X=385640 $Y=935500
X645 354 2 326 1 INV1S $T=388120 920760 1 180 $X=386880 $Y=920380
X646 348 2 330 1 INV1S $T=388740 981240 0 180 $X=387500 $Y=975820
X647 332 2 353 1 INV1S $T=388120 1001400 1 0 $X=388120 $Y=995980
X648 391 2 360 1 INV1S $T=395560 930840 1 180 $X=394320 $Y=930460
X649 369 2 364 1 INV1S $T=394320 1001400 0 0 $X=394320 $Y=1001020
X650 375 2 362 1 INV1S $T=395560 910680 1 0 $X=395560 $Y=905260
X651 383 2 371 1 INV1S $T=398040 940920 1 180 $X=396800 $Y=940540
X652 379 2 363 1 INV1S $T=397420 961080 1 0 $X=397420 $Y=955660
X653 381 2 366 1 INV1S $T=397420 991320 1 0 $X=397420 $Y=985900
X654 382 2 365 1 INV1S $T=399280 961080 0 0 $X=399280 $Y=960700
X655 380 2 376 1 INV1S $T=399280 971160 1 0 $X=399280 $Y=965740
X656 408 2 377 1 INV1S $T=401760 1001400 0 180 $X=400520 $Y=995980
X657 385 2 386 1 INV1S $T=401760 961080 0 0 $X=401760 $Y=960700
X658 395 2 349 1 INV1S $T=402380 900600 0 0 $X=402380 $Y=900220
X659 18 2 401 1 INV1S $T=404240 1041720 1 0 $X=404240 $Y=1036300
X660 405 2 409 1 INV1S $T=405480 1001400 0 0 $X=405480 $Y=1001020
X661 406 2 398 1 INV1S $T=405480 1011480 0 0 $X=405480 $Y=1011100
X662 389 2 413 1 INV1S $T=407340 910680 0 0 $X=407340 $Y=910300
X663 397 2 403 1 INV1S $T=407960 940920 0 0 $X=407960 $Y=940540
X664 411 2 404 1 INV1S $T=407960 971160 1 0 $X=407960 $Y=965740
X665 393 2 414 1 INV1S $T=408580 930840 1 0 $X=408580 $Y=925420
X666 390 2 417 1 INV1S $T=408580 1021560 0 0 $X=408580 $Y=1021180
X667 416 2 394 1 INV1S $T=410440 951000 1 180 $X=409200 $Y=950620
X668 427 2 421 1 INV1S $T=412920 1041720 1 0 $X=412920 $Y=1036300
X669 392 2 432 1 INV1S $T=414160 920760 1 0 $X=414160 $Y=915340
X670 437 2 444 1 INV1S $T=416020 900600 0 0 $X=416020 $Y=900220
X671 450 2 426 1 INV1S $T=417260 1001400 1 180 $X=416020 $Y=1001020
X672 433 2 439 1 INV1S $T=417260 1031640 1 0 $X=417260 $Y=1026220
X673 492 2 445 1 INV1S $T=421600 961080 1 180 $X=420360 $Y=960700
X674 459 2 461 1 INV1S $T=422220 930840 0 0 $X=422220 $Y=930460
X675 463 2 425 1 INV1S $T=423460 951000 1 180 $X=422220 $Y=950620
X676 457 2 458 1 INV1S $T=422220 1011480 0 0 $X=422220 $Y=1011100
X677 464 2 451 1 INV1S $T=423460 1041720 1 180 $X=422220 $Y=1041340
X678 480 2 443 1 INV1S $T=424080 981240 0 180 $X=422840 $Y=975820
X679 472 2 465 1 INV1S $T=425940 991320 0 0 $X=425940 $Y=990940
X680 479 2 454 1 INV1S $T=427800 1011480 1 180 $X=426560 $Y=1011100
X681 486 2 449 1 INV1S $T=428420 920760 1 180 $X=427180 $Y=920380
X682 491 2 483 1 INV1S $T=429660 991320 1 180 $X=428420 $Y=990940
X683 467 2 477 1 INV1S $T=430280 910680 0 0 $X=430280 $Y=910300
X684 489 2 499 1 INV1S $T=430900 930840 0 0 $X=430900 $Y=930460
X685 516 2 505 1 INV1S $T=437100 951000 1 180 $X=435860 $Y=950620
X686 517 2 506 1 INV1S $T=437100 971160 0 180 $X=435860 $Y=965740
X687 539 2 484 1 INV1S $T=437100 1051800 1 180 $X=435860 $Y=1051420
X688 514 2 509 1 INV1S $T=437720 940920 1 0 $X=437720 $Y=935500
X689 522 2 507 1 INV1S $T=438960 1011480 1 180 $X=437720 $Y=1011100
X690 528 2 513 1 INV1S $T=440200 1061880 0 180 $X=438960 $Y=1056460
X691 501 2 529 1 INV1S $T=439580 910680 0 0 $X=439580 $Y=910300
X692 526 2 482 1 INV1S $T=440820 1001400 1 0 $X=440820 $Y=995980
X693 531 2 515 1 INV1S $T=441440 981240 1 0 $X=441440 $Y=975820
X694 551 2 534 1 INV1S $T=445160 951000 0 180 $X=443920 $Y=945580
X695 545 2 512 1 INV1S $T=443920 1031640 1 0 $X=443920 $Y=1026220
X696 31 2 524 1 INV1S $T=447020 900600 1 180 $X=445780 $Y=900220
X697 555 2 530 1 INV1S $T=447640 981240 1 180 $X=446400 $Y=980860
X698 577 2 503 1 INV1S $T=448260 981240 0 180 $X=447020 $Y=975820
X699 561 2 548 1 INV1S $T=448880 951000 1 180 $X=447640 $Y=950620
X700 541 2 564 1 INV1S $T=448260 1001400 0 0 $X=448260 $Y=1001020
X701 567 2 549 1 INV1S $T=450120 1061880 0 180 $X=448880 $Y=1056460
X702 568 2 553 1 INV1S $T=450740 910680 1 180 $X=449500 $Y=910300
X703 579 2 546 1 INV1S $T=453840 1011480 0 0 $X=453840 $Y=1011100
X704 586 2 565 1 INV1S $T=455080 1051800 0 180 $X=453840 $Y=1046380
X705 35 2 544 1 INV1S $T=456320 900600 1 180 $X=455080 $Y=900220
X706 594 2 583 1 INV1S $T=457560 951000 1 180 $X=456320 $Y=950620
X707 595 2 584 1 INV1S $T=457560 971160 1 180 $X=456320 $Y=970780
X708 589 2 573 1 INV1S $T=456320 1021560 1 0 $X=456320 $Y=1016140
X709 590 2 569 1 INV1S $T=457560 1031640 0 180 $X=456320 $Y=1026220
X710 600 2 488 1 INV1S $T=458180 940920 0 180 $X=456940 $Y=935500
X711 596 2 580 1 INV1S $T=458180 981240 1 180 $X=456940 $Y=980860
X712 593 2 624 1 INV1S $T=461280 1021560 1 0 $X=461280 $Y=1016140
X713 614 2 582 1 INV1S $T=461900 930840 0 0 $X=461900 $Y=930460
X714 615 2 606 1 INV1S $T=461900 1001400 1 0 $X=461900 $Y=995980
X715 616 2 602 1 INV1S $T=462520 920760 0 0 $X=462520 $Y=920380
X716 617 2 610 1 INV1S $T=462520 1051800 0 0 $X=462520 $Y=1051420
X717 41 2 39 1 INV1S $T=463760 900600 0 0 $X=463760 $Y=900220
X718 621 2 588 1 INV1S $T=464380 930840 0 0 $X=464380 $Y=930460
X719 599 2 626 1 INV1S $T=464380 1071960 1 0 $X=464380 $Y=1066540
X720 630 2 609 1 INV1S $T=466860 951000 1 180 $X=465620 $Y=950620
X721 625 2 620 1 INV1S $T=465620 1031640 0 0 $X=465620 $Y=1031260
X722 611 2 641 1 INV1S $T=466860 940920 0 0 $X=466860 $Y=940540
X723 633 2 598 1 INV1S $T=468100 971160 1 180 $X=466860 $Y=970780
X724 619 2 628 1 INV1S $T=466860 1011480 1 0 $X=466860 $Y=1006060
X725 639 2 623 1 INV1S $T=468720 981240 1 180 $X=467480 $Y=980860
X726 647 2 634 1 INV1S $T=469340 1041720 0 180 $X=468100 $Y=1036300
X727 655 2 627 1 INV1S $T=470580 910680 0 180 $X=469340 $Y=905260
X728 523 2 649 1 INV1S $T=469340 1011480 1 0 $X=469340 $Y=1006060
X729 652 2 592 1 INV1S $T=471820 1011480 1 0 $X=471820 $Y=1006060
X730 646 2 651 1 INV1S $T=471820 1031640 0 0 $X=471820 $Y=1031260
X731 674 2 648 1 INV1S $T=473680 910680 1 180 $X=472440 $Y=910300
X732 654 2 665 1 INV1S $T=473060 971160 1 0 $X=473060 $Y=965740
X733 669 2 638 1 INV1S $T=474920 1051800 0 180 $X=473680 $Y=1046380
X734 677 2 673 1 INV1S $T=476160 1051800 0 180 $X=474920 $Y=1046380
X735 676 2 645 1 INV1S $T=475540 951000 0 0 $X=475540 $Y=950620
X736 663 2 690 1 INV1S $T=477400 930840 1 0 $X=477400 $Y=925420
X737 689 2 668 1 INV1S $T=478640 991320 0 180 $X=477400 $Y=985900
X738 686 2 669 1 INV1S $T=478640 1051800 0 180 $X=477400 $Y=1046380
X739 669 2 684 1 INV1S $T=477400 1061880 1 0 $X=477400 $Y=1056460
X740 649 2 694 1 INV1S $T=478640 1011480 1 0 $X=478640 $Y=1006060
X741 700 2 658 1 INV1S $T=483600 1071960 0 180 $X=482360 $Y=1066540
X742 707 2 664 1 INV1S $T=484220 940920 1 180 $X=482980 $Y=940540
X743 703 2 682 1 INV1S $T=484220 1011480 1 180 $X=482980 $Y=1011100
X744 708 2 693 1 INV1S $T=484220 1031640 1 180 $X=482980 $Y=1031260
X745 711 2 656 1 INV1S $T=484840 1051800 0 180 $X=483600 $Y=1046380
X746 706 2 687 1 INV1S $T=485460 1071960 1 0 $X=485460 $Y=1066540
X747 730 2 691 1 INV1S $T=487940 951000 0 180 $X=486700 $Y=945580
X748 720 2 714 1 INV1S $T=486700 1001400 1 0 $X=486700 $Y=995980
X749 723 2 718 1 INV1S $T=489180 920760 1 0 $X=489180 $Y=915340
X750 728 2 692 1 INV1S $T=489180 971160 1 0 $X=489180 $Y=965740
X751 713 2 699 1 INV1S $T=490420 910680 0 0 $X=490420 $Y=910300
X752 729 2 724 1 INV1S $T=490420 930840 0 0 $X=490420 $Y=930460
X753 736 2 719 1 INV1S $T=491660 961080 0 0 $X=491660 $Y=960700
X754 740 2 721 1 INV1S $T=491660 1051800 0 0 $X=491660 $Y=1051420
X755 742 2 732 1 INV1S $T=492280 981240 0 0 $X=492280 $Y=980860
X756 757 2 739 1 INV1S $T=495380 1011480 0 180 $X=494140 $Y=1006060
X757 762 2 726 1 INV1S $T=496000 1041720 0 180 $X=494760 $Y=1036300
X758 759 2 747 1 INV1S $T=496000 1021560 0 0 $X=496000 $Y=1021180
X759 760 2 749 1 INV1S $T=497240 1071960 0 180 $X=496000 $Y=1066540
X760 784 2 701 1 INV1S $T=498480 951000 0 180 $X=497240 $Y=945580
X761 771 2 763 1 INV1S $T=497860 971160 0 0 $X=497860 $Y=970780
X762 754 2 758 1 INV1S $T=498480 920760 1 0 $X=498480 $Y=915340
X763 765 2 738 1 INV1S $T=498480 940920 0 0 $X=498480 $Y=940540
X764 773 2 735 1 INV1S $T=499100 1031640 0 0 $X=499100 $Y=1031260
X765 781 2 774 1 INV1S $T=502200 961080 1 180 $X=500960 $Y=960700
X766 780 2 772 1 INV1S $T=501580 991320 0 0 $X=501580 $Y=990940
X767 786 2 779 1 INV1S $T=502820 1001400 1 180 $X=501580 $Y=1001020
X768 794 2 745 1 INV1S $T=504060 981240 0 180 $X=502820 $Y=975820
X769 791 2 778 1 INV1S $T=504680 930840 0 180 $X=503440 $Y=925420
X770 798 2 737 1 INV1S $T=504680 1051800 1 180 $X=503440 $Y=1051420
X771 764 2 810 1 INV1S $T=504680 1011480 1 0 $X=504680 $Y=1006060
X772 796 2 804 1 INV1S $T=506540 961080 1 0 $X=506540 $Y=955660
X773 808 2 793 1 INV1S $T=507780 1071960 0 180 $X=506540 $Y=1066540
X774 788 2 807 1 INV1S $T=507780 910680 0 0 $X=507780 $Y=910300
X775 815 2 748 1 INV1S $T=509640 1031640 1 180 $X=508400 $Y=1031260
X776 51 2 816 1 INV1S $T=508400 1071960 0 0 $X=508400 $Y=1071580
X777 824 2 767 1 INV1S $T=510260 930840 0 0 $X=510260 $Y=930460
X778 821 2 802 1 INV1S $T=510260 1031640 0 0 $X=510260 $Y=1031260
X779 846 2 825 1 INV1S $T=513360 1061880 0 180 $X=512120 $Y=1056460
X780 831 2 803 1 INV1S $T=514600 961080 0 180 $X=513360 $Y=955660
X781 834 2 789 1 INV1S $T=515840 971160 1 180 $X=514600 $Y=970780
X782 845 2 814 1 INV1S $T=516460 920760 1 180 $X=515220 $Y=920380
X783 850 2 837 1 INV1S $T=518320 1051800 1 180 $X=517080 $Y=1051420
X784 848 2 836 1 INV1S $T=518940 991320 1 180 $X=517700 $Y=990940
X785 857 2 838 1 INV1S $T=520800 1031640 1 180 $X=519560 $Y=1031260
X786 858 2 841 1 INV1S $T=520800 1011480 1 0 $X=520800 $Y=1006060
X787 859 2 854 1 INV1S $T=523280 1071960 0 180 $X=522040 $Y=1066540
X788 869 2 826 1 INV1S $T=523900 910680 0 0 $X=523900 $Y=910300
X789 882 2 835 1 INV1S $T=525140 971160 0 180 $X=523900 $Y=965740
X790 872 2 878 1 INV1S $T=523900 1011480 1 0 $X=523900 $Y=1006060
X791 879 2 870 1 INV1S $T=526380 951000 1 180 $X=525140 $Y=950620
X792 886 2 881 1 INV1S $T=528860 1041720 1 180 $X=527620 $Y=1041340
X793 893 2 877 1 INV1S $T=529480 981240 1 180 $X=528240 $Y=980860
X794 887 2 865 1 INV1S $T=528860 951000 1 0 $X=528860 $Y=945580
X795 890 2 867 1 INV1S $T=530100 971160 1 180 $X=528860 $Y=970780
X796 884 2 905 1 INV1S $T=529480 930840 0 0 $X=529480 $Y=930460
X797 929 2 847 1 INV1S $T=532580 951000 1 180 $X=531340 $Y=950620
X798 906 2 888 1 INV1S $T=532580 1071960 0 180 $X=531340 $Y=1066540
X799 902 2 873 1 INV1S $T=532580 1051800 0 0 $X=532580 $Y=1051420
X800 897 2 885 1 INV1S $T=535060 910680 0 0 $X=535060 $Y=910300
X801 925 2 916 1 INV1S $T=536300 991320 0 180 $X=535060 $Y=985900
X802 927 2 895 1 INV1S $T=536300 1051800 1 180 $X=535060 $Y=1051420
X803 934 2 914 1 INV1S $T=536920 1041720 0 180 $X=535680 $Y=1036300
X804 928 2 909 1 INV1S $T=537540 1001400 1 180 $X=536300 $Y=1001020
X805 958 2 908 1 INV1S $T=541260 920760 1 180 $X=540020 $Y=920380
X806 913 2 941 1 INV1S $T=540020 1051800 1 0 $X=540020 $Y=1046380
X807 948 2 901 1 INV1S $T=542500 1021560 1 180 $X=541260 $Y=1021180
X808 945 2 926 1 INV1S $T=543120 910680 1 180 $X=541880 $Y=910300
X809 970 2 932 1 INV1S $T=543740 971160 0 180 $X=542500 $Y=965740
X810 959 2 933 1 INV1S $T=544980 1021560 1 180 $X=543740 $Y=1021180
X811 954 2 949 1 INV1S $T=545600 961080 1 180 $X=544360 $Y=960700
X812 962 2 946 1 INV1S $T=546840 1051800 1 180 $X=545600 $Y=1051420
X813 985 2 950 1 INV1S $T=548080 1001400 1 180 $X=546840 $Y=1001020
X814 982 2 952 1 INV1S $T=550560 930840 1 180 $X=549320 $Y=930460
X815 957 2 921 1 INV1S $T=549320 971160 0 0 $X=549320 $Y=970780
X816 979 2 978 1 INV1S $T=549940 981240 0 0 $X=549940 $Y=980860
X817 984 2 953 1 INV1S $T=551800 1041720 1 180 $X=550560 $Y=1041340
X818 983 2 992 1 INV1S $T=553040 961080 0 0 $X=553040 $Y=960700
X819 991 2 980 1 INV1S $T=553040 1021560 1 0 $X=553040 $Y=1016140
X820 996 2 972 1 INV1S $T=554280 1051800 0 180 $X=553040 $Y=1046380
X821 1010 2 987 1 INV1S $T=556140 940920 0 180 $X=554900 $Y=935500
X822 1001 2 966 1 INV1S $T=556760 910680 1 180 $X=555520 $Y=910300
X823 1024 2 999 1 INV1S $T=558000 1041720 0 180 $X=556760 $Y=1036300
X824 1018 2 1009 1 INV1S $T=558000 1061880 1 180 $X=556760 $Y=1061500
X825 1014 2 998 1 INV1S $T=558620 981240 0 180 $X=557380 $Y=975820
X826 1005 2 939 1 INV1S $T=558000 961080 1 0 $X=558000 $Y=955660
X827 1023 2 1008 1 INV1S $T=560480 1021560 1 180 $X=559240 $Y=1021180
X828 1020 2 981 1 INV1S $T=559240 1071960 1 0 $X=559240 $Y=1066540
X829 1030 2 1002 1 INV1S $T=561100 920760 1 180 $X=559860 $Y=920380
X830 1053 2 1011 1 INV1S $T=561720 1001400 0 180 $X=560480 $Y=995980
X831 1034 2 1003 1 INV1S $T=562960 930840 1 180 $X=561720 $Y=930460
X832 1057 2 1029 1 INV1S $T=564820 961080 1 180 $X=563580 $Y=960700
X833 1040 2 1022 1 INV1S $T=564820 951000 1 0 $X=564820 $Y=945580
X834 994 2 1048 1 INV1S $T=566060 1021560 1 0 $X=566060 $Y=1016140
X835 1056 2 1052 1 INV1S $T=567920 1061880 0 0 $X=567920 $Y=1061500
X836 1063 2 1050 1 INV1S $T=569780 920760 0 180 $X=568540 $Y=915340
X837 1068 2 1038 1 INV1S $T=571020 940920 1 0 $X=571020 $Y=935500
X838 1047 2 1066 1 INV1S $T=572260 1001400 0 180 $X=571020 $Y=995980
X839 1062 2 1028 1 INV1S $T=572880 900600 0 0 $X=572880 $Y=900220
X840 1055 2 1083 1 INV1S $T=572880 951000 0 0 $X=572880 $Y=950620
X841 1088 2 1060 1 INV1S $T=574740 940920 0 180 $X=573500 $Y=935500
X842 1086 2 1051 1 INV1S $T=574740 1031640 0 180 $X=573500 $Y=1026220
X843 1094 2 1073 1 INV1S $T=575360 1041720 1 180 $X=574120 $Y=1041340
X844 1097 2 1080 1 INV1S $T=576600 981240 1 180 $X=575360 $Y=980860
X845 1096 2 1085 1 INV1S $T=577220 920760 1 180 $X=575980 $Y=920380
X846 1090 2 1100 1 INV1S $T=577840 991320 0 0 $X=577840 $Y=990940
X847 1112 2 1093 1 INV1S $T=579080 1071960 0 180 $X=577840 $Y=1066540
X848 1116 2 1067 1 INV1S $T=580320 951000 0 180 $X=579080 $Y=945580
X849 1107 2 1081 1 INV1S $T=580940 1011480 1 180 $X=579700 $Y=1011100
X850 1133 2 1092 1 INV1S $T=581560 1021560 0 180 $X=580320 $Y=1016140
X851 1124 2 1109 1 INV1S $T=582180 900600 1 180 $X=580940 $Y=900220
X852 1064 2 1118 1 INV1S $T=580940 961080 0 0 $X=580940 $Y=960700
X853 1143 2 1101 1 INV1S $T=582180 1041720 0 180 $X=580940 $Y=1036300
X854 1111 2 1121 1 INV1S $T=580940 1051800 0 0 $X=580940 $Y=1051420
X855 1131 2 1110 1 INV1S $T=583420 1011480 1 180 $X=582180 $Y=1011100
X856 1125 2 1113 1 INV1S $T=582800 910680 0 0 $X=582800 $Y=910300
X857 1126 2 1089 1 INV1S $T=582800 971160 0 0 $X=582800 $Y=970780
X858 1137 2 1139 1 INV1S $T=586520 1051800 0 0 $X=586520 $Y=1051420
X859 1159 2 1102 1 INV1S $T=588380 1071960 0 180 $X=587140 $Y=1066540
X860 1141 2 1134 1 INV1S $T=587760 940920 0 0 $X=587760 $Y=940540
X861 1146 2 1129 1 INV1S $T=589620 920760 1 180 $X=588380 $Y=920380
X862 1163 2 1132 1 INV1S $T=589620 991320 0 180 $X=588380 $Y=985900
X863 1155 2 1106 1 INV1S $T=591480 1031640 1 180 $X=590240 $Y=1031260
X864 1161 2 1114 1 INV1S $T=592720 930840 0 0 $X=592720 $Y=930460
X865 1166 2 1157 1 INV1S $T=593960 971160 1 180 $X=592720 $Y=970780
X866 1171 2 1160 1 INV1S $T=594580 1071960 0 180 $X=593340 $Y=1066540
X867 72 2 69 1 INV1S $T=594580 900600 0 0 $X=594580 $Y=900220
X868 1158 2 1192 1 INV1S $T=594580 1031640 0 0 $X=594580 $Y=1031260
X869 1186 2 1154 1 INV1S $T=597060 1011480 1 180 $X=595820 $Y=1011100
X870 1190 2 1168 1 INV1S $T=598920 1001400 1 180 $X=597680 $Y=1001020
X871 1173 2 1151 1 INV1S $T=598300 910680 1 0 $X=598300 $Y=905260
X872 75 2 1128 1 INV1S $T=599540 940920 1 180 $X=598300 $Y=940540
X873 1189 2 1147 1 INV1S $T=598300 961080 0 0 $X=598300 $Y=960700
X874 1199 2 1178 1 INV1S $T=600780 1051800 0 180 $X=599540 $Y=1046380
X875 1196 2 1177 1 INV1S $T=600160 940920 0 0 $X=600160 $Y=940540
X876 1194 2 1214 1 INV1S $T=602020 951000 0 0 $X=602020 $Y=950620
X877 1145 2 1201 1 INV1S $T=602020 971160 0 0 $X=602020 $Y=970780
X878 1202 2 1209 1 INV1S $T=603880 1041720 1 0 $X=603880 $Y=1036300
X879 1224 2 70 1 INV1S $T=606360 910680 0 180 $X=605120 $Y=905260
X880 1221 2 1181 1 INV1S $T=606360 920760 0 180 $X=605120 $Y=915340
X881 1183 2 1227 1 INV1S $T=605120 1051800 0 0 $X=605120 $Y=1051420
X882 1268 2 1215 1 INV1S $T=606980 1011480 1 180 $X=605740 $Y=1011100
X883 1223 2 1176 1 INV1S $T=606360 920760 0 0 $X=606360 $Y=920380
X884 1218 2 1211 1 INV1S $T=606360 991320 1 0 $X=606360 $Y=985900
X885 1233 2 1182 1 INV1S $T=608220 961080 1 180 $X=606980 $Y=960700
X886 1234 2 1195 1 INV1S $T=608840 971160 1 180 $X=607600 $Y=970780
X887 1228 2 1212 1 INV1S $T=608840 1071960 1 0 $X=608840 $Y=1066540
X888 1236 2 1208 1 INV1S $T=610080 1011480 1 0 $X=610080 $Y=1006060
X889 1251 2 1238 1 INV1S $T=612560 1031640 0 180 $X=611320 $Y=1026220
X890 1256 2 81 1 INV1S $T=613180 930840 1 180 $X=611940 $Y=930460
X891 1219 2 1247 1 INV1S $T=611940 1001400 1 0 $X=611940 $Y=995980
X892 1248 2 1198 1 INV1S $T=613180 1021560 0 0 $X=613180 $Y=1021180
X893 1271 2 1254 1 INV1S $T=616280 961080 0 180 $X=615040 $Y=955660
X894 1265 2 82 1 INV1S $T=616900 910680 0 180 $X=615660 $Y=905260
X895 1292 2 1249 1 INV1S $T=616900 1051800 1 180 $X=615660 $Y=1051420
X896 1274 2 1252 1 INV1S $T=617520 981240 1 180 $X=616280 $Y=980860
X897 1267 2 1243 1 INV1S $T=618140 920760 1 180 $X=616900 $Y=920380
X898 1262 2 1232 1 INV1S $T=617520 940920 0 0 $X=617520 $Y=940540
X899 1286 2 1244 1 INV1S $T=619380 1041720 1 180 $X=618140 $Y=1041340
X900 1276 2 1255 1 INV1S $T=620000 971160 1 180 $X=618760 $Y=970780
X901 1272 2 83 1 INV1S $T=619380 920760 0 0 $X=619380 $Y=920380
X902 1253 2 1277 1 INV1S $T=619380 1031640 1 0 $X=619380 $Y=1026220
X903 1273 2 1281 1 INV1S $T=620000 1011480 1 0 $X=620000 $Y=1006060
X904 1285 2 88 1 INV1S $T=621240 920760 1 0 $X=621240 $Y=915340
X905 1308 2 1280 1 INV1S $T=623720 940920 1 180 $X=622480 $Y=940540
X906 1309 2 1278 1 INV1S $T=626820 961080 1 180 $X=625580 $Y=960700
X907 1306 2 1291 1 INV1S $T=626820 1021560 0 180 $X=625580 $Y=1016140
X908 1319 2 1293 1 INV1S $T=628060 930840 1 180 $X=626820 $Y=930460
X909 1310 2 1295 1 INV1S $T=627440 991320 0 0 $X=627440 $Y=990940
X910 1312 2 1294 1 INV1S $T=628060 991320 1 0 $X=628060 $Y=985900
X911 1290 2 1307 1 INV1S $T=629300 1041720 1 180 $X=628060 $Y=1041340
X912 1317 2 1311 1 INV1S $T=628680 1061880 1 0 $X=628680 $Y=1056460
X913 1302 2 1314 1 INV1S $T=630540 1031640 0 180 $X=629300 $Y=1026220
X914 43 2 1305 1 INV1S $T=632400 930840 1 180 $X=631160 $Y=930460
X915 1342 2 1332 1 INV1S $T=635500 981240 0 180 $X=634260 $Y=975820
X916 43 2 1237 1 INV1S $T=635500 991320 0 180 $X=634260 $Y=985900
X917 1343 2 1325 1 INV1S $T=635500 1021560 0 180 $X=634260 $Y=1016140
X918 1348 2 1337 1 INV1S $T=636740 940920 0 180 $X=635500 $Y=935500
X919 1341 2 1299 1 INV1S $T=636120 910680 0 0 $X=636120 $Y=910300
X920 43 2 1344 1 INV1S $T=637360 1021560 1 0 $X=637360 $Y=1016140
X921 1356 2 1289 1 INV1S $T=639220 920760 1 180 $X=637980 $Y=920380
X922 1326 2 1353 1 INV1S $T=637980 1061880 0 0 $X=637980 $Y=1061500
X923 1333 2 1339 1 INV1S $T=637980 1071960 1 0 $X=637980 $Y=1066540
X924 1346 2 1328 1 INV1S $T=638600 951000 1 0 $X=638600 $Y=945580
X925 1359 2 96 1 INV1S $T=639840 900600 0 0 $X=639840 $Y=900220
X926 1365 2 1338 1 INV1S $T=641080 1031640 0 180 $X=639840 $Y=1026220
X927 1367 2 1324 1 INV1S $T=642320 991320 0 180 $X=641080 $Y=985900
X928 1368 2 1347 1 INV1S $T=642320 1011480 0 180 $X=641080 $Y=1006060
X929 1382 2 1363 1 INV1S $T=642940 1041720 1 180 $X=641700 $Y=1041340
X930 1362 2 98 1 INV1S $T=642940 920760 1 0 $X=642940 $Y=915340
X931 1396 2 1357 1 INV1S $T=644800 981240 1 180 $X=643560 $Y=980860
X932 1371 2 1381 1 INV1S $T=644180 1001400 1 0 $X=644180 $Y=995980
X933 1331 2 1383 1 INV1S $T=644800 961080 1 0 $X=644800 $Y=955660
X934 1392 2 1369 1 INV1S $T=646660 940920 0 180 $X=645420 $Y=935500
X935 1400 2 1366 1 INV1S $T=648520 951000 0 180 $X=647280 $Y=945580
X936 1370 2 1387 1 INV1S $T=647900 991320 0 0 $X=647900 $Y=990940
X937 1391 2 1398 1 INV1S $T=647900 1041720 0 0 $X=647900 $Y=1041340
X938 1401 2 1394 1 INV1S $T=650380 1031640 1 0 $X=650380 $Y=1026220
X939 1380 2 1358 1 INV1S $T=651000 961080 0 0 $X=651000 $Y=960700
X940 1445 2 1377 1 INV1S $T=652860 1011480 1 180 $X=651620 $Y=1011100
X941 1410 2 1264 1 INV1S $T=652860 1021560 1 180 $X=651620 $Y=1021180
X942 1421 2 1404 1 INV1S $T=653480 991320 1 180 $X=652240 $Y=990940
X943 1430 2 1412 1 INV1S $T=656580 920760 1 180 $X=655340 $Y=920380
X944 1419 2 100 1 INV1S $T=655340 940920 1 0 $X=655340 $Y=935500
X945 1388 2 1437 1 INV1S $T=655340 1051800 0 0 $X=655340 $Y=1051420
X946 1418 2 95 1 INV1S $T=655960 910680 1 0 $X=655960 $Y=905260
X947 1433 2 101 1 INV1S $T=657200 920760 0 180 $X=655960 $Y=915340
X948 1452 2 1397 1 INV1S $T=657200 961080 0 180 $X=655960 $Y=955660
X949 1436 2 1415 1 INV1S $T=657820 951000 0 180 $X=656580 $Y=945580
X950 75 2 1420 1 INV1S $T=658440 940920 0 0 $X=658440 $Y=940540
X951 1435 2 1386 1 INV1S $T=659060 1071960 1 0 $X=659060 $Y=1066540
X952 1468 2 1444 1 INV1S $T=662160 1001400 0 180 $X=660920 $Y=995980
X953 1446 2 1440 1 INV1S $T=662160 1031640 1 0 $X=662160 $Y=1026220
X954 1458 2 1457 1 INV1S $T=663400 1061880 1 0 $X=663400 $Y=1056460
X955 1461 2 106 1 INV1S $T=664020 920760 0 0 $X=664020 $Y=920380
X956 1453 2 1406 1 INV1S $T=665260 971160 1 0 $X=665260 $Y=965740
X957 1469 2 1414 1 INV1S $T=666500 991320 0 180 $X=665260 $Y=985900
X958 1476 2 110 1 INV1S $T=667740 920760 1 180 $X=666500 $Y=920380
X959 1478 2 1467 1 INV1S $T=668980 981240 1 180 $X=667740 $Y=980860
X960 1470 2 1425 1 INV1S $T=667740 1001400 1 0 $X=667740 $Y=995980
X961 1479 2 109 1 INV1S $T=668980 1051800 1 180 $X=667740 $Y=1051420
X962 1483 2 1462 1 INV1S $T=669600 940920 0 180 $X=668360 $Y=935500
X963 1472 2 1385 1 INV1S $T=668360 1061880 0 0 $X=668360 $Y=1061500
X964 1495 2 1482 1 INV1S $T=672080 951000 0 180 $X=670840 $Y=945580
X965 1504 2 1413 1 INV1S $T=672700 961080 0 180 $X=671460 $Y=955660
X966 1494 2 1487 1 INV1S $T=673320 1011480 0 180 $X=672080 $Y=1006060
X967 114 2 1474 1 INV1S $T=673320 1071960 0 0 $X=673320 $Y=1071580
X968 1502 2 1475 1 INV1S $T=675180 971160 0 180 $X=673940 $Y=965740
X969 1491 2 1473 1 INV1S $T=673940 1021560 1 0 $X=673940 $Y=1016140
X970 1506 2 1455 1 INV1S $T=675800 1041720 0 0 $X=675800 $Y=1041340
X971 1481 2 119 1 INV1S $T=677040 910680 1 0 $X=677040 $Y=905260
X972 1510 2 1519 1 INV1S $T=677660 1021560 1 0 $X=677660 $Y=1016140
X973 1523 2 117 1 INV1S $T=680140 920760 1 180 $X=678900 $Y=920380
X974 1514 2 1520 1 INV1S $T=680760 1031640 1 0 $X=680760 $Y=1026220
X975 1530 2 1488 1 INV1S $T=680760 1061880 1 0 $X=680760 $Y=1056460
X976 1542 2 1498 1 INV1S $T=682620 940920 1 180 $X=681380 $Y=940540
X977 1526 2 1521 1 INV1S $T=681380 981240 1 0 $X=681380 $Y=975820
X978 1541 2 1529 1 INV1S $T=684480 971160 0 180 $X=683240 $Y=965740
X979 1544 2 1490 1 INV1S $T=684480 1031640 0 180 $X=683240 $Y=1026220
X980 1540 2 1464 1 INV1S $T=683860 1071960 0 0 $X=683860 $Y=1071580
X981 1509 2 1545 1 INV1S $T=685100 961080 1 0 $X=685100 $Y=955660
X982 1547 2 122 1 INV1S $T=685720 930840 0 0 $X=685720 $Y=930460
X983 1531 2 1558 1 INV1S $T=686960 1021560 0 0 $X=686960 $Y=1021180
X984 1565 2 1522 1 INV1S $T=688820 920760 0 180 $X=687580 $Y=915340
X985 1570 2 1512 1 INV1S $T=688820 930840 1 180 $X=687580 $Y=930460
X986 1563 2 1492 1 INV1S $T=689440 1051800 0 180 $X=688200 $Y=1046380
X987 1568 2 1538 1 INV1S $T=690060 981240 1 180 $X=688820 $Y=980860
X988 1571 2 1518 1 INV1S $T=690680 961080 0 180 $X=689440 $Y=955660
X989 1572 2 1505 1 INV1S $T=690680 981240 0 180 $X=689440 $Y=975820
X990 1564 2 1569 1 INV1S $T=689440 1011480 1 0 $X=689440 $Y=1006060
X991 1576 2 1539 1 INV1S $T=691920 1001400 0 0 $X=691920 $Y=1001020
X992 1555 2 1573 1 INV1S $T=693160 1031640 1 0 $X=693160 $Y=1026220
X993 1560 2 1537 1 INV1S $T=693780 951000 1 0 $X=693780 $Y=945580
X994 1586 2 1554 1 INV1S $T=693780 981240 0 0 $X=693780 $Y=980860
X995 43 2 1578 1 INV1S $T=695020 1051800 1 180 $X=693780 $Y=1051420
X996 1598 2 1588 1 INV1S $T=697500 940920 0 180 $X=696260 $Y=935500
X997 1612 2 1546 1 INV1S $T=698740 1051800 0 180 $X=697500 $Y=1046380
X998 1599 2 1557 1 INV1S $T=698740 940920 0 0 $X=698740 $Y=940540
X999 1608 2 1595 1 INV1S $T=699980 930840 1 0 $X=699980 $Y=925420
X1000 133 2 1587 1 INV1S $T=702460 900600 1 180 $X=701220 $Y=900220
X1001 1622 2 1607 1 INV1S $T=702460 910680 1 180 $X=701220 $Y=910300
X1002 1620 2 1561 1 INV1S $T=701840 971160 1 0 $X=701840 $Y=965740
X1003 1638 2 1577 1 INV1S $T=703080 1051800 1 180 $X=701840 $Y=1051420
X1004 1616 2 1615 1 INV1S $T=703080 1071960 1 0 $X=703080 $Y=1066540
X1005 1631 2 1589 1 INV1S $T=703700 1001400 0 0 $X=703700 $Y=1001020
X1006 1639 2 1543 1 INV1S $T=705560 1021560 1 180 $X=704320 $Y=1021180
X1007 135 2 1636 1 INV1S $T=706180 900600 1 180 $X=704940 $Y=900220
X1008 1609 2 1613 1 INV1S $T=705560 1001400 1 0 $X=705560 $Y=995980
X1009 1642 2 1532 1 INV1S $T=706800 1071960 0 180 $X=705560 $Y=1066540
X1010 1640 2 1597 1 INV1S $T=706180 1011480 1 0 $X=706180 $Y=1006060
X1011 1644 2 1619 1 INV1S $T=706800 1021560 0 0 $X=706800 $Y=1021180
X1012 1646 2 1610 1 INV1S $T=708040 1031640 1 180 $X=706800 $Y=1031260
X1013 1660 2 1652 1 INV1S $T=710520 910680 1 180 $X=709280 $Y=910300
X1014 1664 2 1593 1 INV1S $T=710520 1051800 0 180 $X=709280 $Y=1046380
X1015 1655 2 1614 1 INV1S $T=710520 1061880 0 180 $X=709280 $Y=1056460
X1016 1670 2 1618 1 INV1S $T=711760 951000 0 180 $X=710520 $Y=945580
X1017 1662 2 1667 1 INV1S $T=710520 971160 0 0 $X=710520 $Y=970780
X1018 1674 2 1641 1 INV1S $T=713620 1051800 0 180 $X=712380 $Y=1046380
X1019 1675 2 1637 1 INV1S $T=714240 981240 1 180 $X=713000 $Y=980860
X1020 1673 2 1683 1 INV1S $T=713000 1071960 0 0 $X=713000 $Y=1071580
X1021 1677 2 1661 1 INV1S $T=714240 930840 0 0 $X=714240 $Y=930460
X1022 1650 2 1686 1 INV1S $T=714240 961080 0 0 $X=714240 $Y=960700
X1023 1687 2 1643 1 INV1S $T=718580 920760 0 180 $X=717340 $Y=915340
X1024 1700 2 1645 1 INV1S $T=719200 951000 1 0 $X=719200 $Y=945580
X1025 1680 2 1696 1 INV1S $T=719820 981240 0 0 $X=719820 $Y=980860
X1026 1705 2 1681 1 INV1S $T=721060 991320 0 180 $X=719820 $Y=985900
X1027 1709 2 1634 1 INV1S $T=721060 1031640 1 180 $X=719820 $Y=1031260
X1028 1740 2 1676 1 INV1S $T=721680 1001400 0 180 $X=720440 $Y=995980
X1029 1716 2 1669 1 INV1S $T=722300 1031640 0 180 $X=721060 $Y=1026220
X1030 1684 2 1708 1 INV1S $T=721680 930840 0 0 $X=721680 $Y=930460
X1031 1725 2 1679 1 INV1S $T=726020 930840 1 180 $X=724780 $Y=930460
X1032 1748 2 1690 1 INV1S $T=727260 1031640 1 180 $X=726020 $Y=1031260
X1033 1727 2 1653 1 INV1S $T=727260 971160 1 0 $X=727260 $Y=965740
X1034 1739 2 1651 1 INV1S $T=729120 961080 1 180 $X=727880 $Y=960700
X1035 1745 2 140 1 INV1S $T=729740 951000 0 180 $X=728500 $Y=945580
X1036 1752 2 1697 1 INV1S $T=729740 1011480 1 180 $X=728500 $Y=1011100
X1037 1731 2 1672 1 INV1S $T=728500 1041720 0 0 $X=728500 $Y=1041340
X1038 1735 2 1712 1 INV1S $T=730360 920760 0 180 $X=729120 $Y=915340
X1039 146 2 1730 1 INV1S $T=731600 1071960 0 0 $X=731600 $Y=1071580
X1040 1743 2 1724 1 INV1S $T=732220 1011480 1 0 $X=732220 $Y=1006060
X1041 1753 2 1689 1 INV1S $T=733460 951000 1 0 $X=733460 $Y=945580
X1042 1754 2 1763 1 INV1S $T=734080 1031640 0 0 $X=734080 $Y=1031260
X1043 1757 2 1704 1 INV1S $T=734700 940920 1 0 $X=734700 $Y=935500
X1044 1747 2 1737 1 INV1S $T=735940 1011480 0 180 $X=734700 $Y=1006060
X1045 1749 2 1701 1 INV1S $T=734700 1051800 0 0 $X=734700 $Y=1051420
X1046 1758 2 1726 1 INV1S $T=735940 951000 0 0 $X=735940 $Y=950620
X1047 1764 2 1698 1 INV1S $T=736560 1031640 1 0 $X=736560 $Y=1026220
X1048 1768 2 1746 1 INV1S $T=738420 920760 0 180 $X=737180 $Y=915340
X1049 1772 2 1777 1 INV1S $T=737800 1061880 1 0 $X=737800 $Y=1056460
X1050 1761 2 1760 1 INV1S $T=738420 971160 1 0 $X=738420 $Y=965740
X1051 1775 2 1781 1 INV1S $T=739660 910680 0 0 $X=739660 $Y=910300
X1052 1798 2 1733 1 INV1S $T=743380 1031640 0 180 $X=742140 $Y=1026220
X1053 149 2 1796 1 INV1S $T=744620 981240 1 180 $X=743380 $Y=980860
X1054 1790 2 1786 1 INV1S $T=743380 1051800 1 0 $X=743380 $Y=1046380
X1055 1742 2 1729 1 INV1S $T=744000 961080 0 0 $X=744000 $Y=960700
X1056 1801 2 1774 1 INV1S $T=745240 991320 1 180 $X=744000 $Y=990940
X1057 1802 2 1778 1 INV1S $T=746480 1001400 0 180 $X=745240 $Y=995980
X1058 1792 2 1776 1 INV1S $T=745240 1011480 0 0 $X=745240 $Y=1011100
X1059 1821 2 1815 1 INV1S $T=749580 930840 1 0 $X=749580 $Y=925420
X1060 1813 2 1816 1 INV1S $T=750200 971160 0 0 $X=750200 $Y=970780
X1061 161 2 1784 1 INV1S $T=750200 1071960 0 0 $X=750200 $Y=1071580
X1062 1800 2 1822 1 INV1S $T=750820 1031640 0 0 $X=750820 $Y=1031260
X1063 158 2 1808 1 INV1S $T=751440 910680 0 0 $X=751440 $Y=910300
X1064 163 2 162 1 INV1S $T=753300 900600 1 180 $X=752060 $Y=900220
X1065 1835 2 1793 1 INV1S $T=753300 1061880 1 180 $X=752060 $Y=1061500
X1066 1833 2 1825 1 INV1S $T=753300 1021560 1 0 $X=753300 $Y=1016140
X1067 1832 2 1765 1 INV1S $T=753920 920760 1 0 $X=753920 $Y=915340
X1068 1843 2 1783 1 INV1S $T=756400 940920 0 180 $X=755160 $Y=935500
X1069 1850 2 1823 1 INV1S $T=757020 1061880 1 180 $X=755780 $Y=1061500
X1070 1851 2 1848 1 INV1S $T=758880 940920 0 180 $X=757640 $Y=935500
X1071 1853 2 1828 1 INV1S $T=757640 1001400 1 0 $X=757640 $Y=995980
X1072 1854 2 1819 1 INV1S $T=758260 1041720 0 0 $X=758260 $Y=1041340
X1073 1841 2 1855 1 INV1S $T=758880 1061880 0 0 $X=758880 $Y=1061500
X1074 1862 2 1826 1 INV1S $T=760740 961080 1 180 $X=759500 $Y=960700
X1075 1856 2 1872 1 INV1S $T=760120 981240 0 0 $X=760120 $Y=980860
X1076 1863 2 1846 1 INV1S $T=761980 1041720 1 180 $X=760740 $Y=1041340
X1077 1845 2 1849 1 INV1S $T=761360 1001400 0 0 $X=761360 $Y=1001020
X1078 1866 2 1824 1 INV1S $T=761980 910680 0 0 $X=761980 $Y=910300
X1079 1844 2 1852 1 INV1S $T=763840 961080 1 0 $X=763840 $Y=955660
X1080 1884 2 1847 1 INV1S $T=764460 1031640 1 0 $X=764460 $Y=1026220
X1081 1877 2 1804 1 INV1S $T=765700 951000 1 0 $X=765700 $Y=945580
X1082 1886 2 1860 1 INV1S $T=765700 971160 1 0 $X=765700 $Y=965740
X1083 1874 2 168 1 INV1S $T=766940 910680 0 0 $X=766940 $Y=910300
X1084 1876 2 1869 1 INV1S $T=767560 1031640 1 0 $X=767560 $Y=1026220
X1085 144 2 1908 1 INV1S $T=768180 910680 0 0 $X=768180 $Y=910300
X1086 1896 2 1842 1 INV1S $T=769420 971160 0 180 $X=768180 $Y=965740
X1087 1897 2 1868 1 INV1S $T=768180 991320 0 0 $X=768180 $Y=990940
X1088 1901 2 1889 1 INV1S $T=768800 1001400 0 0 $X=768800 $Y=1001020
X1089 1904 2 1887 1 INV1S $T=770040 1071960 1 180 $X=768800 $Y=1071580
X1090 1879 2 1882 1 INV1S $T=769420 930840 1 0 $X=769420 $Y=925420
X1091 1918 2 1919 1 INV1S $T=771900 1021560 1 0 $X=771900 $Y=1016140
X1092 1928 2 1880 1 INV1S $T=773760 940920 0 180 $X=772520 $Y=935500
X1093 174 2 1814 1 INV1S $T=775000 1071960 1 180 $X=773760 $Y=1071580
X1094 1920 2 1883 1 INV1S $T=774380 1021560 0 0 $X=774380 $Y=1021180
X1095 1903 2 1907 1 INV1S $T=774380 1061880 0 0 $X=774380 $Y=1061500
X1096 1943 2 1932 1 INV1S $T=778100 940920 0 180 $X=776860 $Y=935500
X1097 1946 2 1890 1 INV1S $T=779960 1041720 0 180 $X=778720 $Y=1036300
X1098 1952 2 1936 1 INV1S $T=781200 900600 1 180 $X=779960 $Y=900220
X1099 1934 2 1938 1 INV1S $T=781820 1011480 0 180 $X=780580 $Y=1006060
X1100 176 2 178 1 INV1S $T=781820 900600 0 0 $X=781820 $Y=900220
X1101 1961 2 1924 1 INV1S $T=783060 920760 0 180 $X=781820 $Y=915340
X1102 1953 2 1922 1 INV1S $T=781820 951000 1 0 $X=781820 $Y=945580
X1103 1949 2 1931 1 INV1S $T=782440 1041720 1 0 $X=782440 $Y=1036300
X1104 1959 2 1962 1 INV1S $T=783680 1001400 1 0 $X=783680 $Y=995980
X1105 1958 2 1972 1 INV1S $T=784300 981240 0 0 $X=784300 $Y=980860
X1106 1967 2 1957 1 INV1S $T=785540 1061880 0 180 $X=784300 $Y=1056460
X1107 1937 2 1982 1 INV1S $T=786160 961080 0 0 $X=786160 $Y=960700
X1108 1987 2 1941 1 INV1S $T=789260 1021560 0 180 $X=788020 $Y=1016140
X1109 1975 2 1954 1 INV1S $T=788640 981240 1 0 $X=788640 $Y=975820
X1110 1998 2 1977 1 INV1S $T=792360 910680 1 180 $X=791120 $Y=910300
X1111 2005 2 1965 1 INV1S $T=792980 930840 1 0 $X=792980 $Y=925420
X1112 1999 2 1945 1 INV1S $T=792980 940920 1 0 $X=792980 $Y=935500
X1113 2014 2 1993 1 INV1S $T=794840 1031640 1 180 $X=793600 $Y=1031260
X1114 2018 2 1992 1 INV1S $T=795460 1001400 0 180 $X=794220 $Y=995980
X1115 2010 2 2009 1 INV1S $T=794840 981240 1 0 $X=794840 $Y=975820
X1116 1915 2 2015 1 INV1S $T=795460 930840 1 0 $X=795460 $Y=925420
X1117 2015 2 2013 1 INV1S $T=797320 940920 0 180 $X=796080 $Y=935500
X1118 2027 2 1976 1 INV1S $T=797940 1071960 0 180 $X=796700 $Y=1066540
X1119 2017 2 2024 1 INV1S $T=797320 1021560 1 0 $X=797320 $Y=1016140
X1120 2015 2 2000 1 INV1S $T=797940 930840 1 0 $X=797940 $Y=925420
X1121 2036 2 1914 1 INV1S $T=800420 951000 1 180 $X=799180 $Y=950620
X1122 2045 2 1970 1 INV1S $T=801040 1021560 0 180 $X=799800 $Y=1016140
X1123 2029 2 1991 1 INV1S $T=800420 951000 1 0 $X=800420 $Y=945580
X1124 2031 2 2008 1 INV1S $T=800420 1061880 0 0 $X=800420 $Y=1061500
X1125 2047 2 2023 1 INV1S $T=802900 930840 0 180 $X=801660 $Y=925420
X1126 2040 2 1973 1 INV1S $T=802900 1011480 1 180 $X=801660 $Y=1011100
X1127 2044 2 2028 1 INV1S $T=802900 1041720 1 180 $X=801660 $Y=1041340
X1128 2069 2 2039 1 INV1S $T=804140 981240 1 180 $X=802900 $Y=980860
X1129 2043 2 2016 1 INV1S $T=802900 991320 1 0 $X=802900 $Y=985900
X1130 2059 2 1859 1 INV1S $T=804760 910680 1 180 $X=803520 $Y=910300
X1131 2048 2 2041 1 INV1S $T=804140 1031640 0 0 $X=804140 $Y=1031260
X1132 2083 2 2055 1 INV1S $T=809720 951000 1 180 $X=808480 $Y=950620
X1133 2070 2 2052 1 INV1S $T=809100 1001400 0 0 $X=809100 $Y=1001020
X1134 2081 2 2053 1 INV1S $T=813440 930840 0 180 $X=812200 $Y=925420
X1135 2068 2 1906 1 INV1S $T=812200 940920 0 0 $X=812200 $Y=940540
X1136 2085 2 2087 1 INV1S $T=813440 971160 0 0 $X=813440 $Y=970780
X1137 2092 2 2011 1 INV1S $T=815920 1021560 0 180 $X=814680 $Y=1016140
X1138 2103 2 2086 1 INV1S $T=818400 1011480 1 180 $X=817160 $Y=1011100
X1139 2109 2 2062 1 INV1S $T=818400 1041720 1 180 $X=817160 $Y=1041340
X1140 2095 2 2106 1 INV1S $T=819020 1001400 0 0 $X=819020 $Y=1001020
X1141 2102 2 2096 1 INV1S $T=819640 961080 1 0 $X=819640 $Y=955660
X1142 2119 2 2073 1 INV1S $T=822120 1041720 0 180 $X=820880 $Y=1036300
X1143 2107 2 2104 1 INV1S $T=821500 981240 0 0 $X=821500 $Y=980860
X1144 2118 2 2098 1 INV1S $T=822740 1031640 0 180 $X=821500 $Y=1026220
X1145 2105 2 1974 1 INV1S $T=821500 1051800 0 0 $X=821500 $Y=1051420
X1146 2115 2 2093 1 INV1S $T=823360 940920 0 180 $X=822120 $Y=935500
X1147 2128 2 2117 1 INV1S $T=830180 981240 1 180 $X=828940 $Y=980860
X1148 2123 2 2091 1 INV1S $T=831420 971160 0 180 $X=830180 $Y=965740
X1149 2124 2 2072 1 INV1S $T=832660 1011480 0 0 $X=832660 $Y=1011100
X1150 2131 2 2122 1 INV1S $T=836380 1001400 1 180 $X=835140 $Y=1001020
X1151 2130 2 2114 1 INV1S $T=836380 1011480 1 180 $X=835140 $Y=1011100
X1152 211 2 2125 1 INV1S $T=840100 900600 1 180 $X=838860 $Y=900220
X1153 2132 2 2133 1 INV1S $T=841960 910680 0 0 $X=841960 $Y=910300
X1154 2164 2 2147 1 INV1S $T=865520 930840 1 180 $X=864280 $Y=930460
X1155 210 2 2150 1 INV1S $T=868000 930840 0 180 $X=866760 $Y=925420
X1156 203 2 2175 1 INV1S $T=872960 930840 1 0 $X=872960 $Y=925420
X1157 2166 2 2173 1 INV1S $T=874820 910680 0 180 $X=873580 $Y=905260
X1158 235 2 2176 1 INV1S $T=877300 940920 1 0 $X=877300 $Y=935500
X1159 212 2 2186 1 INV1S $T=881640 920760 1 0 $X=881640 $Y=915340
X1160 2193 2 2198 1 INV1S $T=886600 900600 0 0 $X=886600 $Y=900220
X1161 2199 2 2195 1 INV1S $T=889080 920760 0 180 $X=887840 $Y=915340
X1162 2203 2 2206 1 INV1S $T=893420 940920 1 0 $X=893420 $Y=935500
X1163 2212 2 2211 1 INV1S $T=895900 930840 0 180 $X=894660 $Y=925420
X1164 246 2 2207 1 INV1S $T=898380 930840 0 180 $X=897140 $Y=925420
X1165 246 2 245 1 INV1S $T=897760 910680 1 0 $X=897760 $Y=905260
X1166 246 2 2217 1 INV1S $T=898380 930840 1 0 $X=898380 $Y=925420
X1167 2215 2 2218 1 INV1S $T=900240 920760 1 0 $X=900240 $Y=915340
X1168 247 2 2228 1 INV1S $T=902720 900600 0 0 $X=902720 $Y=900220
X1169 2224 2 2231 1 INV1S $T=904580 920760 0 0 $X=904580 $Y=920380
X1170 2209 2 2236 1 INV1S $T=907060 951000 1 180 $X=905820 $Y=950620
X1171 250 2 2229 1 INV1S $T=906440 920760 0 0 $X=906440 $Y=920380
X1172 252 2 2246 1 INV1S $T=911400 910680 1 0 $X=911400 $Y=905260
X1173 2244 2 2259 1 INV1S $T=920080 951000 1 0 $X=920080 $Y=945580
X1174 2245 2 2260 1 INV1S $T=921320 920760 1 0 $X=921320 $Y=915340
X1175 2247 2 2261 1 INV1S $T=923800 940920 0 0 $X=923800 $Y=940540
X1176 2265 2 2270 1 INV1S $T=927520 930840 1 0 $X=927520 $Y=925420
X1177 2256 2 2272 1 INV1S $T=928760 930840 0 0 $X=928760 $Y=930460
X1178 2276 2 2271 1 INV1S $T=932480 920760 1 0 $X=932480 $Y=915340
X1179 2264 2 2292 1 INV1S $T=941160 940920 1 0 $X=941160 $Y=935500
X1180 2204 2 2294 1 INV1S $T=943640 940920 1 0 $X=943640 $Y=935500
X1181 2170 2 2295 1 INV1S $T=949840 930840 0 180 $X=948600 $Y=925420
X1182 2240 2 2302 1 INV1S $T=960380 951000 0 180 $X=959140 $Y=945580
X1183 273 2 2314 1 INV1S $T=965340 910680 1 0 $X=965340 $Y=905260
X1184 302 305 298 300 2 1 MXL2HS $T=368280 930840 0 180 $X=362700 $Y=925420
X1185 301 7 304 9 2 1 MXL2HS $T=363320 910680 1 0 $X=363320 $Y=905260
X1186 307 305 299 302 2 1 MXL2HS $T=368900 940920 0 180 $X=363320 $Y=935500
X1187 300 308 306 301 2 1 MXL2HS $T=371380 920760 0 180 $X=365800 $Y=915340
X1188 311 318 312 307 2 1 MXL2HS $T=375100 961080 0 180 $X=369520 $Y=955660
X1189 320 318 315 311 2 1 MXL2HS $T=375720 971160 0 180 $X=370140 $Y=965740
X1190 322 318 319 327 2 1 MXL2HS $T=376340 961080 1 0 $X=376340 $Y=955660
X1191 330 318 321 322 2 1 MXL2HS $T=382540 971160 0 180 $X=376960 $Y=965740
X1192 325 308 309 13 2 1 MXL2HS $T=383780 910680 0 180 $X=378200 $Y=905260
X1193 336 308 328 325 2 1 MXL2HS $T=385020 920760 0 180 $X=379440 $Y=915340
X1194 341 305 316 326 2 1 MXL2HS $T=385640 930840 1 180 $X=380060 $Y=930460
X1195 327 329 317 341 2 1 MXL2HS $T=380060 940920 0 0 $X=380060 $Y=940540
X1196 349 11 342 17 2 1 MXL2HS $T=389360 900600 1 180 $X=383780 $Y=900220
X1197 353 358 352 330 2 1 MXL2HS $T=391840 991320 0 180 $X=386260 $Y=985900
X1198 362 11 351 349 2 1 MXL2HS $T=392460 910680 0 180 $X=386880 $Y=905260
X1199 326 308 357 362 2 1 MXL2HS $T=386880 920760 1 0 $X=386880 $Y=915340
X1200 360 305 355 336 2 1 MXL2HS $T=392460 930840 1 180 $X=386880 $Y=930460
X1201 364 358 333 353 2 1 MXL2HS $T=393080 1001400 1 180 $X=387500 $Y=1001020
X1202 371 305 359 360 2 1 MXL2HS $T=395560 940920 1 180 $X=389980 $Y=940540
X1203 363 329 344 371 2 1 MXL2HS $T=390600 951000 1 0 $X=390600 $Y=945580
X1204 365 370 345 363 2 1 MXL2HS $T=396180 961080 0 180 $X=390600 $Y=955660
X1205 376 373 346 365 2 1 MXL2HS $T=397420 971160 0 180 $X=391840 $Y=965740
X1206 377 358 368 366 2 1 MXL2HS $T=397420 991320 0 180 $X=391840 $Y=985900
X1207 366 373 347 386 2 1 MXL2HS $T=395560 981240 1 0 $X=395560 $Y=975820
X1208 398 358 374 377 2 1 MXL2HS $T=403620 1001400 1 180 $X=398040 $Y=1001020
X1209 394 329 387 403 2 1 MXL2HS $T=401140 940920 0 0 $X=401140 $Y=940540
X1210 404 373 384 320 2 1 MXL2HS $T=406720 971160 0 180 $X=401140 $Y=965740
X1211 386 329 402 394 2 1 MXL2HS $T=402380 951000 0 0 $X=402380 $Y=950620
X1212 403 305 410 414 2 1 MXL2HS $T=404860 930840 0 0 $X=404860 $Y=930460
X1213 421 418 396 409 2 1 MXL2HS $T=412920 1041720 0 180 $X=407340 $Y=1036300
X1214 426 358 412 364 2 1 MXL2HS $T=413540 1001400 1 180 $X=407960 $Y=1001020
X1215 417 418 415 398 2 1 MXL2HS $T=413540 1011480 1 180 $X=407960 $Y=1011100
X1216 432 428 420 413 2 1 MXL2HS $T=415400 910680 1 180 $X=409820 $Y=910300
X1217 409 358 431 436 2 1 MXL2HS $T=410440 991320 0 0 $X=410440 $Y=990940
X1218 425 370 429 438 2 1 MXL2HS $T=411680 951000 0 0 $X=411680 $Y=950620
X1219 439 418 399 417 2 1 MXL2HS $T=417260 1021560 1 180 $X=411680 $Y=1021180
X1220 443 373 430 376 2 1 MXL2HS $T=417880 971160 1 180 $X=412300 $Y=970780
X1221 445 370 434 425 2 1 MXL2HS $T=418500 961080 0 180 $X=412920 $Y=955660
X1222 446 370 435 404 2 1 MXL2HS $T=418500 971160 0 180 $X=412920 $Y=965740
X1223 413 428 422 444 2 1 MXL2HS $T=414160 910680 1 0 $X=414160 $Y=905260
X1224 414 428 423 449 2 1 MXL2HS $T=414160 920760 0 0 $X=414160 $Y=920380
X1225 451 418 442 421 2 1 MXL2HS $T=420360 1041720 0 180 $X=414780 $Y=1036300
X1226 436 440 388 445 2 1 MXL2HS $T=415400 981240 0 0 $X=415400 $Y=980860
X1227 454 418 441 426 2 1 MXL2HS $T=420980 1011480 1 180 $X=415400 $Y=1011100
X1228 444 23 400 24 2 1 MXL2HS $T=417880 900600 0 0 $X=417880 $Y=900220
X1229 438 452 424 461 2 1 MXL2HS $T=418500 940920 1 0 $X=418500 $Y=935500
X1230 461 428 447 432 2 1 MXL2HS $T=425940 920760 1 180 $X=420360 $Y=920380
X1231 468 418 456 458 2 1 MXL2HS $T=426560 1021560 1 180 $X=420980 $Y=1021180
X1232 449 428 455 477 2 1 MXL2HS $T=422220 910680 0 0 $X=422220 $Y=910300
X1233 465 440 448 443 2 1 MXL2HS $T=427800 981240 1 180 $X=422220 $Y=980860
X1234 482 466 469 465 2 1 MXL2HS $T=429040 1001400 0 180 $X=423460 $Y=995980
X1235 458 466 474 483 2 1 MXL2HS $T=423460 1001400 0 0 $X=423460 $Y=1001020
X1236 484 481 471 468 2 1 MXL2HS $T=429660 1051800 0 180 $X=424080 $Y=1046380
X1237 485 481 476 451 2 1 MXL2HS $T=430280 1041720 1 180 $X=424700 $Y=1041340
X1238 29 25 27 26 2 1 MXL2HS $T=431520 900600 1 180 $X=425940 $Y=900220
X1239 503 440 490 446 2 1 MXL2HS $T=434000 981240 0 180 $X=428420 $Y=975820
X1240 505 452 478 488 2 1 MXL2HS $T=434620 951000 1 180 $X=429040 $Y=950620
X1241 483 440 498 506 2 1 MXL2HS $T=429660 981240 0 0 $X=429660 $Y=980860
X1242 507 475 487 454 2 1 MXL2HS $T=435240 1011480 1 180 $X=429660 $Y=1011100
X1243 509 452 473 499 2 1 MXL2HS $T=436480 940920 0 180 $X=430900 $Y=935500
X1244 477 25 508 29 2 1 MXL2HS $T=431520 900600 0 0 $X=431520 $Y=900220
X1245 513 481 495 484 2 1 MXL2HS $T=437720 1061880 0 180 $X=432140 $Y=1056460
X1246 506 519 502 505 2 1 MXL2HS $T=440200 961080 0 180 $X=434620 $Y=955660
X1247 515 440 497 503 2 1 MXL2HS $T=440200 981240 0 180 $X=434620 $Y=975820
X1248 530 440 511 515 2 1 MXL2HS $T=442060 981240 1 180 $X=436480 $Y=980860
X1249 524 25 30 544 2 1 MXL2HS $T=439580 900600 0 0 $X=439580 $Y=900220
X1250 534 452 518 509 2 1 MXL2HS $T=445160 940920 0 180 $X=439580 $Y=935500
X1251 529 521 537 524 2 1 MXL2HS $T=440200 910680 1 0 $X=440200 $Y=905260
X1252 546 475 533 507 2 1 MXL2HS $T=445780 1011480 1 180 $X=440200 $Y=1011100
X1253 548 519 538 534 2 1 MXL2HS $T=447020 951000 1 180 $X=441440 $Y=950620
X1254 549 481 540 513 2 1 MXL2HS $T=447020 1061880 0 180 $X=441440 $Y=1056460
X1255 553 521 542 529 2 1 MXL2HS $T=447640 910680 1 180 $X=442060 $Y=910300
X1256 554 466 500 482 2 1 MXL2HS $T=447640 1001400 0 180 $X=442060 $Y=995980
X1257 499 550 527 543 2 1 MXL2HS $T=448880 930840 0 180 $X=443300 $Y=925420
X1258 543 550 494 553 2 1 MXL2HS $T=445160 920760 0 0 $X=445160 $Y=920380
X1259 565 481 558 485 2 1 MXL2HS $T=451360 1051800 0 180 $X=445780 $Y=1046380
X1260 569 481 552 512 2 1 MXL2HS $T=451980 1031640 0 180 $X=446400 $Y=1026220
X1261 573 475 547 546 2 1 MXL2HS $T=452600 1011480 1 180 $X=447020 $Y=1011100
X1262 564 466 562 554 2 1 MXL2HS $T=453220 1001400 0 180 $X=447640 $Y=995980
X1263 544 521 32 33 2 1 MXL2HS $T=448260 900600 0 0 $X=448260 $Y=900220
X1264 580 578 559 530 2 1 MXL2HS $T=455080 981240 1 180 $X=449500 $Y=980860
X1265 488 560 566 582 2 1 MXL2HS $T=450120 940920 1 0 $X=450120 $Y=935500
X1266 583 519 556 548 2 1 MXL2HS $T=455700 951000 1 180 $X=450120 $Y=950620
X1267 584 519 557 572 2 1 MXL2HS $T=456320 961080 1 180 $X=450740 $Y=960700
X1268 598 578 587 584 2 1 MXL2HS $T=460040 981240 0 180 $X=454460 $Y=975820
X1269 582 560 570 602 2 1 MXL2HS $T=455080 930840 0 0 $X=455080 $Y=930460
X1270 602 521 574 588 2 1 MXL2HS $T=461280 920760 1 180 $X=455700 $Y=920380
X1271 606 578 571 564 2 1 MXL2HS $T=461280 1001400 0 180 $X=455700 $Y=995980
X1272 572 519 603 609 2 1 MXL2HS $T=456320 961080 0 0 $X=456320 $Y=960700
X1273 610 605 575 565 2 1 MXL2HS $T=461900 1051800 0 180 $X=456320 $Y=1046380
X1274 33 36 38 39 2 1 MXL2HS $T=456940 900600 0 0 $X=456940 $Y=900220
X1275 592 591 604 606 2 1 MXL2HS $T=456940 1011480 1 0 $X=456940 $Y=1006060
X1276 609 519 607 583 2 1 MXL2HS $T=464380 951000 1 180 $X=458800 $Y=950620
X1277 620 605 581 569 2 1 MXL2HS $T=464380 1031640 1 180 $X=458800 $Y=1031260
X1278 623 578 612 580 2 1 MXL2HS $T=465000 981240 1 180 $X=459420 $Y=980860
X1279 627 36 618 40 2 1 MXL2HS $T=466860 910680 0 180 $X=461280 $Y=905260
X1280 634 638 613 626 2 1 MXL2HS $T=469960 1051800 0 180 $X=464380 $Y=1046380
X1281 626 638 629 549 2 1 MXL2HS $T=469960 1061880 0 180 $X=464380 $Y=1056460
X1282 628 578 635 645 2 1 MXL2HS $T=465000 1001400 1 0 $X=465000 $Y=995980
X1283 648 521 631 627 2 1 MXL2HS $T=471200 910680 1 180 $X=465620 $Y=910300
X1284 588 521 640 648 2 1 MXL2HS $T=465620 920760 0 0 $X=465620 $Y=920380
X1285 624 591 636 628 2 1 MXL2HS $T=465620 1021560 1 0 $X=465620 $Y=1016140
X1286 651 605 637 624 2 1 MXL2HS $T=471820 1031640 0 180 $X=466240 $Y=1026220
X1287 656 638 644 610 2 1 MXL2HS $T=473060 1051800 1 180 $X=467480 $Y=1051420
X1288 645 650 632 641 2 1 MXL2HS $T=474300 951000 1 180 $X=468720 $Y=950620
X1289 641 650 653 664 2 1 MXL2HS $T=469340 940920 0 0 $X=469340 $Y=940540
X1290 665 659 608 598 2 1 MXL2HS $T=474920 971160 1 180 $X=469340 $Y=970780
X1291 668 659 642 623 2 1 MXL2HS $T=475540 981240 1 180 $X=469960 $Y=980860
X1292 673 605 657 651 2 1 MXL2HS $T=476160 1041720 0 180 $X=470580 $Y=1036300
X1293 658 638 671 673 2 1 MXL2HS $T=471820 1061880 1 0 $X=471820 $Y=1056460
X1294 682 591 660 573 2 1 MXL2HS $T=478640 1011480 1 180 $X=473060 $Y=1011100
X1295 687 684 662 658 2 1 MXL2HS $T=479880 1071960 0 180 $X=474300 $Y=1066540
X1296 692 659 681 665 2 1 MXL2HS $T=481120 971160 0 180 $X=475540 $Y=965740
X1297 693 686 667 620 2 1 MXL2HS $T=481120 1031640 1 180 $X=475540 $Y=1031260
X1298 664 650 666 691 2 1 MXL2HS $T=476160 940920 0 0 $X=476160 $Y=940540
X1299 695 659 678 668 2 1 MXL2HS $T=481740 981240 1 180 $X=476160 $Y=980860
X1300 691 650 685 701 2 1 MXL2HS $T=479260 951000 1 0 $X=479260 $Y=945580
X1301 714 675 679 682 2 1 MXL2HS $T=486700 1011480 0 180 $X=481120 $Y=1006060
X1302 718 715 680 699 2 1 MXL2HS $T=487940 920760 0 180 $X=482360 $Y=915340
X1303 719 659 688 692 2 1 MXL2HS $T=487940 971160 0 180 $X=482360 $Y=965740
X1304 726 686 710 634 2 1 MXL2HS $T=489180 1041720 0 180 $X=483600 $Y=1036300
X1305 735 686 722 693 2 1 MXL2HS $T=491040 1031640 1 180 $X=485460 $Y=1031260
X1306 737 684 725 721 2 1 MXL2HS $T=491660 1051800 0 180 $X=486080 $Y=1046380
X1307 721 684 698 656 2 1 MXL2HS $T=491660 1051800 1 180 $X=486080 $Y=1051420
X1308 690 715 716 718 2 1 MXL2HS $T=492280 920760 1 180 $X=486700 $Y=920380
X1309 724 715 683 690 2 1 MXL2HS $T=492280 930840 0 180 $X=486700 $Y=925420
X1310 738 715 717 724 2 1 MXL2HS $T=492280 940920 0 180 $X=486700 $Y=935500
X1311 739 675 727 592 2 1 MXL2HS $T=492900 1011480 0 180 $X=487320 $Y=1006060
X1312 747 686 709 726 2 1 MXL2HS $T=494140 1021560 1 180 $X=488560 $Y=1021180
X1313 749 684 712 687 2 1 MXL2HS $T=494140 1071960 0 180 $X=488560 $Y=1066540
X1314 701 650 743 738 2 1 MXL2HS $T=489800 951000 1 0 $X=489800 $Y=945580
X1315 699 715 752 758 2 1 MXL2HS $T=491660 920760 1 0 $X=491660 $Y=915340
X1316 745 744 755 763 2 1 MXL2HS $T=492280 971160 0 0 $X=492280 $Y=970780
X1317 748 686 756 735 2 1 MXL2HS $T=492280 1031640 0 0 $X=492280 $Y=1031260
X1318 763 744 734 719 2 1 MXL2HS $T=499100 971160 0 180 $X=493520 $Y=965740
X1319 772 768 731 714 2 1 MXL2HS $T=499720 991320 1 180 $X=494140 $Y=990940
X1320 774 744 741 732 2 1 MXL2HS $T=500340 961080 1 180 $X=494760 $Y=960700
X1321 778 753 761 767 2 1 MXL2HS $T=502200 930840 0 180 $X=496620 $Y=925420
X1322 779 675 751 739 2 1 MXL2HS $T=502200 1011480 0 180 $X=496620 $Y=1006060
X1323 758 753 776 778 2 1 MXL2HS $T=497240 920760 0 0 $X=497240 $Y=920380
X1324 789 783 777 745 2 1 MXL2HS $T=504680 971160 1 180 $X=499100 $Y=970780
X1325 793 787 766 749 2 1 MXL2HS $T=505300 1071960 0 180 $X=499720 $Y=1066540
X1326 801 797 769 747 2 1 MXL2HS $T=507160 1021560 1 180 $X=501580 $Y=1021180
X1327 802 797 770 748 2 1 MXL2HS $T=507160 1031640 1 180 $X=501580 $Y=1031260
X1328 803 799 790 774 2 1 MXL2HS $T=507780 961080 1 180 $X=502200 $Y=960700
X1329 805 768 785 772 2 1 MXL2HS $T=508400 991320 1 180 $X=502820 $Y=990940
X1330 810 768 800 779 2 1 MXL2HS $T=509640 1001400 1 180 $X=504060 $Y=1001020
X1331 767 753 775 814 2 1 MXL2HS $T=504680 930840 1 0 $X=504680 $Y=925420
X1332 825 819 806 737 2 1 MXL2HS $T=511500 1051800 1 180 $X=505920 $Y=1051420
X1333 826 560 809 50 2 1 MXL2HS $T=512120 920760 0 180 $X=506540 $Y=915340
X1334 814 753 812 807 2 1 MXL2HS $T=512740 920760 1 180 $X=507160 $Y=920380
X1335 804 799 817 803 2 1 MXL2HS $T=513360 961080 0 180 $X=507780 $Y=955660
X1336 807 753 828 54 2 1 MXL2HS $T=509020 910680 0 0 $X=509020 $Y=910300
X1337 816 787 52 793 2 1 MXL2HS $T=514600 1071960 0 180 $X=509020 $Y=1066540
X1338 835 783 829 789 2 1 MXL2HS $T=517080 971160 0 180 $X=511500 $Y=965740
X1339 837 819 813 825 2 1 MXL2HS $T=517080 1051800 1 180 $X=511500 $Y=1051420
X1340 838 797 822 801 2 1 MXL2HS $T=517700 1031640 1 180 $X=512120 $Y=1031260
X1341 841 53 820 810 2 1 MXL2HS $T=518320 1001400 1 180 $X=512740 $Y=1001020
X1342 854 787 823 816 2 1 MXL2HS $T=520800 1071960 0 180 $X=515220 $Y=1066540
X1343 865 860 842 847 2 1 MXL2HS $T=523280 951000 0 180 $X=517700 $Y=945580
X1344 867 799 852 804 2 1 MXL2HS $T=523900 971160 0 180 $X=518320 $Y=965740
X1345 873 819 861 837 2 1 MXL2HS $T=525140 1051800 1 180 $X=519560 $Y=1051420
X1346 877 768 853 836 2 1 MXL2HS $T=526380 981240 1 180 $X=520800 $Y=980860
X1347 870 799 833 835 2 1 MXL2HS $T=527000 961080 1 180 $X=521420 $Y=960700
X1348 881 797 863 838 2 1 MXL2HS $T=527620 1031640 1 180 $X=522040 $Y=1031260
X1349 878 862 866 841 2 1 MXL2HS $T=528240 1001400 1 180 $X=522660 $Y=1001020
X1350 847 860 875 870 2 1 MXL2HS $T=528860 951000 0 180 $X=523280 $Y=945580
X1351 885 840 849 826 2 1 MXL2HS $T=529480 920760 0 180 $X=523900 $Y=915340
X1352 888 787 864 854 2 1 MXL2HS $T=530100 1071960 0 180 $X=524520 $Y=1066540
X1353 895 819 876 873 2 1 MXL2HS $T=531340 1051800 1 180 $X=525760 $Y=1051420
X1354 909 862 883 878 2 1 MXL2HS $T=534440 1001400 1 180 $X=528860 $Y=1001020
X1355 914 912 896 881 2 1 MXL2HS $T=535680 1041720 1 180 $X=530100 $Y=1041340
X1356 915 860 898 865 2 1 MXL2HS $T=536300 951000 0 180 $X=530720 $Y=945580
X1357 916 911 899 877 2 1 MXL2HS $T=536300 981240 1 180 $X=530720 $Y=980860
X1358 921 911 907 867 2 1 MXL2HS $T=536920 971160 1 180 $X=531340 $Y=970780
X1359 908 840 918 926 2 1 MXL2HS $T=532580 920760 0 0 $X=532580 $Y=920380
X1360 904 840 851 908 2 1 MXL2HS $T=533200 930840 1 0 $X=533200 $Y=925420
X1361 905 924 839 904 2 1 MXL2HS $T=538780 930840 1 180 $X=533200 $Y=930460
X1362 930 787 920 888 2 1 MXL2HS $T=539400 1071960 0 180 $X=533820 $Y=1066540
X1363 932 799 922 916 2 1 MXL2HS $T=540020 971160 0 180 $X=534440 $Y=965740
X1364 933 912 923 901 2 1 MXL2HS $T=540020 1021560 1 180 $X=534440 $Y=1021180
X1365 926 840 903 60 2 1 MXL2HS $T=541880 910680 1 180 $X=536300 $Y=910300
X1366 946 941 919 895 2 1 MXL2HS $T=543740 1051800 1 180 $X=538160 $Y=1051420
X1367 949 860 910 932 2 1 MXL2HS $T=544360 961080 1 180 $X=538780 $Y=960700
X1368 950 862 937 909 2 1 MXL2HS $T=544360 1001400 1 180 $X=538780 $Y=1001020
X1369 952 924 936 905 2 1 MXL2HS $T=544980 930840 1 180 $X=539400 $Y=930460
X1370 953 912 938 914 2 1 MXL2HS $T=544980 1041720 1 180 $X=539400 $Y=1041340
X1371 966 840 956 885 2 1 MXL2HS $T=548700 910680 1 180 $X=543120 $Y=910300
X1372 969 862 947 950 2 1 MXL2HS $T=549320 1001400 0 180 $X=543740 $Y=995980
X1373 972 941 964 946 2 1 MXL2HS $T=550560 1051800 0 180 $X=544980 $Y=1046380
X1374 977 860 961 949 2 1 MXL2HS $T=551180 961080 1 180 $X=545600 $Y=960700
X1375 978 911 951 921 2 1 MXL2HS $T=551180 981240 0 180 $X=545600 $Y=975820
X1376 980 912 944 933 2 1 MXL2HS $T=551800 1021560 1 180 $X=546220 $Y=1021180
X1377 998 911 990 978 2 1 MXL2HS $T=556760 981240 0 180 $X=551180 $Y=975820
X1378 1002 997 986 987 2 1 MXL2HS $T=557380 920760 1 180 $X=551800 $Y=920380
X1379 1003 997 989 952 2 1 MXL2HS $T=557380 930840 1 180 $X=551800 $Y=930460
X1380 999 971 974 953 2 1 MXL2HS $T=557380 1041720 1 180 $X=551800 $Y=1041340
X1381 1008 971 973 980 2 1 MXL2HS $T=558000 1021560 1 180 $X=552420 $Y=1021180
X1382 1009 943 975 981 2 1 MXL2HS $T=558000 1071960 0 180 $X=552420 $Y=1066540
X1383 1028 65 1015 966 2 1 MXL2HS $T=562340 900600 1 180 $X=556760 $Y=900220
X1384 1031 1007 993 1011 2 1 MXL2HS $T=562960 1001400 1 180 $X=557380 $Y=1001020
X1385 1032 971 1000 972 2 1 MXL2HS $T=563580 1041720 1 180 $X=558000 $Y=1041340
X1386 1038 997 1021 1022 2 1 MXL2HS $T=564820 951000 0 180 $X=559240 $Y=945580
X1387 1035 943 1025 1009 2 1 MXL2HS $T=564820 1061880 1 180 $X=559240 $Y=1061500
X1388 1022 992 1006 1029 2 1 MXL2HS $T=566060 961080 0 180 $X=560480 $Y=955660
X1389 1046 1042 1019 998 2 1 MXL2HS $T=567300 971160 1 180 $X=561720 $Y=970780
X1390 1048 1007 1036 1008 2 1 MXL2HS $T=567300 1021560 1 180 $X=561720 $Y=1021180
X1391 1050 997 1016 1002 2 1 MXL2HS $T=567920 920760 1 180 $X=562340 $Y=920380
X1392 1051 1007 1037 1032 2 1 MXL2HS $T=567920 1031640 0 180 $X=562340 $Y=1026220
X1393 1052 943 1033 1035 2 1 MXL2HS $T=567920 1071960 0 180 $X=562340 $Y=1066540
X1394 1060 997 1039 1038 2 1 MXL2HS $T=569780 940920 0 180 $X=564200 $Y=935500
X1395 1080 1042 1044 1066 2 1 MXL2HS $T=574120 981240 1 180 $X=568540 $Y=980860
X1396 1081 1077 1054 1048 2 1 MXL2HS $T=574120 1021560 0 180 $X=568540 $Y=1016140
X1397 1067 997 1079 1083 2 1 MXL2HS $T=569160 951000 1 0 $X=569160 $Y=945580
X1398 1066 1077 1072 1031 2 1 MXL2HS $T=574740 1011480 0 180 $X=569160 $Y=1006060
X1399 1085 1082 1043 1060 2 1 MXL2HS $T=575360 920760 1 180 $X=569780 $Y=920380
X1400 1092 1077 1087 1051 2 1 MXL2HS $T=578460 1021560 1 180 $X=572880 $Y=1021180
X1401 1101 971 1091 1073 2 1 MXL2HS $T=579080 1041720 0 180 $X=573500 $Y=1036300
X1402 1109 66 1074 1028 2 1 MXL2HS $T=580320 900600 1 180 $X=574740 $Y=900220
X1403 1110 1077 1095 1092 2 1 MXL2HS $T=580320 1021560 0 180 $X=574740 $Y=1016140
X1404 1113 1082 1075 1050 2 1 MXL2HS $T=580940 920760 0 180 $X=575360 $Y=915340
X1405 1114 1082 1098 1003 2 1 MXL2HS $T=580940 930840 1 180 $X=575360 $Y=930460
X1406 1118 1042 1105 1100 2 1 MXL2HS $T=582180 971160 1 180 $X=576600 $Y=970780
X1407 1121 1108 1059 1102 2 1 MXL2HS $T=582800 1061880 0 180 $X=577220 $Y=1056460
X1408 1100 1042 1119 1080 2 1 MXL2HS $T=577840 981240 0 0 $X=577840 $Y=980860
X1409 1106 1077 1115 1101 2 1 MXL2HS $T=577840 1031640 0 0 $X=577840 $Y=1031260
X1410 1129 1082 1103 1085 2 1 MXL2HS $T=585280 920760 1 180 $X=579700 $Y=920380
X1411 1083 1128 1104 1089 2 1 MXL2HS $T=585900 961080 0 180 $X=580320 $Y=955660
X1412 1102 1108 1123 1093 2 1 MXL2HS $T=585900 1071960 0 180 $X=580320 $Y=1066540
X1413 1132 1042 1122 1110 2 1 MXL2HS $T=586520 991320 0 180 $X=580940 $Y=985900
X1414 1134 1128 1099 1067 2 1 MXL2HS $T=587140 951000 0 180 $X=581560 $Y=945580
X1415 1139 1108 1120 1121 2 1 MXL2HS $T=588380 1061880 0 180 $X=582800 $Y=1056460
X1416 69 68 67 1109 2 1 MXL2HS $T=589000 900600 1 180 $X=583420 $Y=900220
X1417 1147 1128 1135 1132 2 1 MXL2HS $T=590240 961080 1 180 $X=584660 $Y=960700
X1418 1151 1148 1130 1113 2 1 MXL2HS $T=591480 910680 1 180 $X=585900 $Y=910300
X1419 1157 1152 1127 1114 2 1 MXL2HS $T=592720 971160 1 180 $X=587140 $Y=970780
X1420 1154 1162 1138 1081 2 1 MXL2HS $T=594580 1011480 1 180 $X=589000 $Y=1011100
X1421 1160 1108 1136 1139 2 1 MXL2HS $T=594580 1061880 0 180 $X=589000 $Y=1056460
X1422 1168 1162 1140 1154 2 1 MXL2HS $T=595820 1011480 0 180 $X=590240 $Y=1006060
X1423 70 1148 1169 1176 2 1 MXL2HS $T=591480 910680 0 0 $X=591480 $Y=910300
X1424 1177 1170 1144 1134 2 1 MXL2HS $T=597060 940920 1 180 $X=591480 $Y=940540
X1425 1178 1108 1150 1160 2 1 MXL2HS $T=597060 1051800 1 180 $X=591480 $Y=1051420
X1426 1181 1148 1164 1129 2 1 MXL2HS $T=597680 920760 0 180 $X=592100 $Y=915340
X1427 1182 1175 1165 1118 2 1 MXL2HS $T=597680 961080 1 180 $X=592100 $Y=960700
X1428 1192 1188 1179 1106 2 1 MXL2HS $T=600160 1021560 1 180 $X=594580 $Y=1021180
X1429 1195 1152 1184 1157 2 1 MXL2HS $T=600780 971160 1 180 $X=595200 $Y=970780
X1430 1176 1170 1174 1201 2 1 MXL2HS $T=598300 930840 0 0 $X=598300 $Y=930460
X1431 1208 1162 1185 1192 2 1 MXL2HS $T=604500 1011480 1 180 $X=598920 $Y=1011100
X1432 1211 1162 1167 1168 2 1 MXL2HS $T=605120 1001400 0 180 $X=599540 $Y=995980
X1433 1214 1175 1203 1147 2 1 MXL2HS $T=605740 961080 1 180 $X=600160 $Y=960700
X1434 1215 1188 1204 1198 2 1 MXL2HS $T=605740 1021560 0 180 $X=600160 $Y=1016140
X1435 77 1193 1205 1151 2 1 MXL2HS $T=606360 900600 1 180 $X=600780 $Y=900220
X1436 1201 1152 1191 1215 2 1 MXL2HS $T=600780 981240 0 0 $X=600780 $Y=980860
X1437 1209 1210 1153 1227 2 1 MXL2HS $T=602640 1041720 0 0 $X=602640 $Y=1041340
X1438 1212 76 1180 78 2 1 MXL2HS $T=603260 1061880 0 0 $X=603260 $Y=1061500
X1439 1232 1170 1220 1177 2 1 MXL2HS $T=609460 940920 1 180 $X=603880 $Y=940540
X1440 1198 1188 1197 1238 2 1 MXL2HS $T=604500 1031640 1 0 $X=604500 $Y=1026220
X1441 1243 1170 1225 1214 2 1 MXL2HS $T=610700 930840 1 180 $X=605120 $Y=930460
X1442 1244 1210 1226 1178 2 1 MXL2HS $T=610700 1051800 0 180 $X=605120 $Y=1046380
X1443 1238 1210 1206 1209 2 1 MXL2HS $T=612560 1041720 0 180 $X=606980 $Y=1036300
X1444 82 1193 1239 1181 2 1 MXL2HS $T=613180 910680 0 180 $X=607600 $Y=905260
X1445 1227 76 1245 1249 2 1 MXL2HS $T=607600 1051800 0 0 $X=607600 $Y=1051420
X1446 83 1250 1231 1242 2 1 MXL2HS $T=614420 920760 1 180 $X=608840 $Y=920380
X1447 1252 1222 1230 1208 2 1 MXL2HS $T=614420 991320 0 180 $X=608840 $Y=985900
X1448 1249 76 1246 1212 2 1 MXL2HS $T=614420 1061880 1 180 $X=608840 $Y=1061500
X1449 1254 1175 1240 1247 2 1 MXL2HS $T=615660 971160 0 180 $X=610080 $Y=965740
X1450 81 1170 1229 1254 2 1 MXL2HS $T=610700 940920 0 0 $X=610700 $Y=940540
X1451 1255 1175 1241 1211 2 1 MXL2HS $T=616280 971160 1 180 $X=610700 $Y=970780
X1452 1247 1222 1258 1264 2 1 MXL2HS $T=612560 1011480 1 0 $X=612560 $Y=1006060
X1453 1278 1175 1266 1252 2 1 MXL2HS $T=621240 971160 0 180 $X=615660 $Y=965740
X1454 1277 1188 1275 1244 2 1 MXL2HS $T=623100 1041720 0 180 $X=617520 $Y=1036300
X1455 84 1193 1282 1280 2 1 MXL2HS $T=618140 910680 1 0 $X=618140 $Y=905260
X1456 1291 1288 1261 1277 2 1 MXL2HS $T=624340 1021560 0 180 $X=618760 $Y=1016140
X1457 1293 1250 1283 1182 2 1 MXL2HS $T=624960 930840 1 180 $X=619380 $Y=930460
X1458 1242 1279 1216 1294 2 1 MXL2HS $T=619380 961080 1 0 $X=619380 $Y=955660
X1459 1280 1279 1270 1295 2 1 MXL2HS $T=620000 951000 0 0 $X=620000 $Y=950620
X1460 1299 1250 1287 1243 2 1 MXL2HS $T=626200 920760 1 180 $X=620620 $Y=920380
X1461 1294 1222 1263 1281 2 1 MXL2HS $T=626200 991320 1 180 $X=620620 $Y=990940
X1462 1301 1298 1284 1195 2 1 MXL2HS $T=626820 971160 1 180 $X=621240 $Y=970780
X1463 1289 1250 1297 1293 2 1 MXL2HS $T=621860 930840 1 0 $X=621860 $Y=925420
X1464 1281 1288 1304 1307 2 1 MXL2HS $T=623100 1011480 0 0 $X=623100 $Y=1011100
X1465 1307 1322 1316 1311 2 1 MXL2HS $T=632400 1051800 1 180 $X=626820 $Y=1051420
X1466 1325 1288 1315 1314 2 1 MXL2HS $T=633640 1021560 0 180 $X=628060 $Y=1016140
X1467 1328 1279 1303 1278 2 1 MXL2HS $T=634260 961080 0 180 $X=628680 $Y=955660
X1468 1295 1222 1257 1325 2 1 MXL2HS $T=628680 1001400 1 0 $X=628680 $Y=995980
X1469 1314 1188 1327 1335 2 1 MXL2HS $T=629920 1041720 1 0 $X=629920 $Y=1036300
X1470 88 1250 1329 1337 2 1 MXL2HS $T=630540 920760 0 0 $X=630540 $Y=920380
X1471 1311 1322 1269 1339 2 1 MXL2HS $T=630540 1061880 0 0 $X=630540 $Y=1061500
X1472 1337 1279 1318 1324 2 1 MXL2HS $T=636740 951000 0 180 $X=631160 $Y=945580
X1473 1347 1351 1323 1338 2 1 MXL2HS $T=639840 1011480 0 180 $X=634260 $Y=1006060
X1474 1358 1298 1334 1255 2 1 MXL2HS $T=640460 971160 1 180 $X=634880 $Y=970780
X1475 1324 1351 1330 1347 2 1 MXL2HS $T=641700 1001400 0 180 $X=636120 $Y=995980
X1476 1338 1188 1352 1363 2 1 MXL2HS $T=636740 1041720 1 0 $X=636740 $Y=1036300
X1477 1363 1322 1336 1353 2 1 MXL2HS $T=642940 1051800 1 180 $X=637360 $Y=1051420
X1478 95 90 1364 1369 2 1 MXL2HS $T=638600 910680 0 0 $X=638600 $Y=910300
X1479 1369 1361 1354 1357 2 1 MXL2HS $T=644180 940920 0 180 $X=638600 $Y=935500
X1480 1357 1298 1349 1381 2 1 MXL2HS $T=640460 971160 0 0 $X=640460 $Y=970780
X1481 1366 1279 1355 1383 2 1 MXL2HS $T=641080 951000 1 0 $X=641080 $Y=945580
X1482 1353 97 1375 1385 2 1 MXL2HS $T=641080 1061880 0 0 $X=641080 $Y=1061500
X1483 1339 97 1376 1386 2 1 MXL2HS $T=641080 1071960 1 0 $X=641080 $Y=1066540
X1484 98 1361 1378 1366 2 1 MXL2HS $T=641700 930840 1 0 $X=641700 $Y=925420
X1485 1264 1372 1360 1394 2 1 MXL2HS $T=642940 1031640 1 0 $X=642940 $Y=1026220
X1486 1377 1372 1393 1398 2 1 MXL2HS $T=643560 1021560 1 0 $X=643560 $Y=1016140
X1487 1383 1298 1374 1387 2 1 MXL2HS $T=645420 961080 0 0 $X=645420 $Y=960700
X1488 1387 1351 1399 1404 2 1 MXL2HS $T=645420 1001400 1 0 $X=645420 $Y=995980
X1489 1406 1403 1395 1332 2 1 MXL2HS $T=651620 971160 1 180 $X=646040 $Y=970780
X1490 1381 1351 1405 1377 2 1 MXL2HS $T=646660 1011480 1 0 $X=646660 $Y=1006060
X1491 1397 1298 1408 1411 2 1 MXL2HS $T=647280 971160 1 0 $X=647280 $Y=965740
X1492 1412 1361 1402 1232 2 1 MXL2HS $T=653480 930840 0 180 $X=647900 $Y=925420
X1493 100 1361 1373 1413 2 1 MXL2HS $T=648520 940920 1 0 $X=648520 $Y=935500
X1494 101 1361 1389 1415 2 1 MXL2HS $T=649140 920760 1 0 $X=649140 $Y=915340
X1495 1415 1420 1407 1397 2 1 MXL2HS $T=656580 951000 0 180 $X=651000 $Y=945580
X1496 1404 1351 1416 1425 2 1 MXL2HS $T=651000 1001400 1 0 $X=651000 $Y=995980
X1497 1411 1403 1409 1414 2 1 MXL2HS $T=657820 981240 1 180 $X=652240 $Y=980860
X1498 1394 1424 1431 1440 2 1 MXL2HS $T=654100 1031640 1 0 $X=654100 $Y=1026220
X1499 105 1441 104 1299 2 1 MXL2HS $T=660920 900600 1 180 $X=655340 $Y=900220
X1500 1444 1351 1423 1291 2 1 MXL2HS $T=660920 1011480 0 180 $X=655340 $Y=1006060
X1501 106 1441 1422 1412 2 1 MXL2HS $T=663400 920760 1 180 $X=657820 $Y=920380
X1502 1335 1424 1379 1455 2 1 MXL2HS $T=658440 1041720 1 0 $X=658440 $Y=1036300
X1503 1398 1424 1432 1437 2 1 MXL2HS $T=658440 1051800 1 0 $X=658440 $Y=1046380
X1504 1437 1424 1429 1457 2 1 MXL2HS $T=659060 1051800 0 0 $X=659060 $Y=1051420
X1505 108 1441 1447 1289 2 1 MXL2HS $T=665260 910680 1 180 $X=659680 $Y=910300
X1506 1462 1456 1448 1328 2 1 MXL2HS $T=665260 940920 1 180 $X=659680 $Y=940540
X1507 1386 1428 1390 1464 2 1 MXL2HS $T=659680 1071960 0 0 $X=659680 $Y=1071580
X1508 1385 1428 1427 1474 2 1 MXL2HS $T=662780 1071960 1 0 $X=662780 $Y=1066540
X1509 1413 1420 1465 1475 2 1 MXL2HS $T=663400 961080 1 0 $X=663400 $Y=955660
X1510 1482 1420 1459 1358 2 1 MXL2HS $T=670840 940920 1 180 $X=665260 $Y=940540
X1511 1487 1471 1451 1473 2 1 MXL2HS $T=672080 1021560 0 180 $X=666500 $Y=1016140
X1512 1474 1428 112 1488 2 1 MXL2HS $T=666500 1071960 0 0 $X=666500 $Y=1071580
X1513 1440 1471 1485 1490 2 1 MXL2HS $T=667120 1031640 1 0 $X=667120 $Y=1026220
X1514 1455 1424 1466 1492 2 1 MXL2HS $T=667740 1051800 1 0 $X=667740 $Y=1046380
X1515 110 1441 1442 1498 2 1 MXL2HS $T=668980 920760 0 0 $X=668980 $Y=920380
X1516 1457 1428 1497 116 2 1 MXL2HS $T=670220 1061880 0 0 $X=670220 $Y=1061500
X1517 117 1456 1480 1462 2 1 MXL2HS $T=676420 940920 0 180 $X=670840 $Y=935500
X1518 1414 1503 1496 1487 2 1 MXL2HS $T=677040 1001400 0 180 $X=671460 $Y=995980
X1519 115 1441 118 1512 2 1 MXL2HS $T=672700 900600 0 0 $X=672700 $Y=900220
X1520 1498 1456 1501 1518 2 1 MXL2HS $T=673940 940920 0 0 $X=673940 $Y=940540
X1521 1473 1471 1449 1519 2 1 MXL2HS $T=673940 1021560 0 0 $X=673940 $Y=1021180
X1522 1490 1471 1499 1520 2 1 MXL2HS $T=673940 1031640 1 0 $X=673940 $Y=1026220
X1523 1521 1515 1484 1505 2 1 MXL2HS $T=680140 981240 0 180 $X=674560 $Y=975820
X1524 1475 1477 1460 1521 2 1 MXL2HS $T=675800 971160 0 0 $X=675800 $Y=970780
X1525 122 1456 1500 1482 2 1 MXL2HS $T=682000 940920 0 180 $X=676420 $Y=935500
X1526 1529 1477 1508 1406 2 1 MXL2HS $T=682000 971160 0 180 $X=676420 $Y=965740
X1527 1464 120 1493 1532 2 1 MXL2HS $T=677040 1071960 0 0 $X=677040 $Y=1071580
X1528 1522 1441 1533 1537 2 1 MXL2HS $T=678900 920760 1 0 $X=678900 $Y=915340
X1529 1425 1503 1511 1539 2 1 MXL2HS $T=678900 1001400 0 0 $X=678900 $Y=1001020
X1530 1519 1471 1536 1543 2 1 MXL2HS $T=680140 1021560 0 0 $X=680140 $Y=1021180
X1531 1492 1534 1517 1546 2 1 MXL2HS $T=680760 1051800 1 0 $X=680760 $Y=1046380
X1532 119 124 1524 1545 2 1 MXL2HS $T=682000 910680 0 0 $X=682000 $Y=910300
X1533 1505 1515 1548 1538 2 1 MXL2HS $T=682620 981240 1 0 $X=682620 $Y=975820
X1534 1538 1515 1527 1554 2 1 MXL2HS $T=682620 981240 0 0 $X=682620 $Y=980860
X1535 1512 1456 1535 1557 2 1 MXL2HS $T=683240 940920 1 0 $X=683240 $Y=935500
X1536 109 1534 1528 1558 2 1 MXL2HS $T=683240 1051800 0 0 $X=683240 $Y=1051420
X1537 125 124 1551 1522 2 1 MXL2HS $T=683860 910680 1 0 $X=683860 $Y=905260
X1538 1545 1477 1552 1561 2 1 MXL2HS $T=684480 971160 1 0 $X=684480 $Y=965740
X1539 1562 1477 1549 1467 2 1 MXL2HS $T=690060 971160 1 180 $X=684480 $Y=970780
X1540 1539 1503 1525 1569 2 1 MXL2HS $T=685100 1001400 0 0 $X=685100 $Y=1001020
X1541 1520 1553 1559 1573 2 1 MXL2HS $T=685720 1031640 1 0 $X=685720 $Y=1026220
X1542 1488 1556 1566 1577 2 1 MXL2HS $T=686340 1061880 1 0 $X=686340 $Y=1056460
X1543 1587 124 128 96 2 1 MXL2HS $T=695640 910680 1 180 $X=690060 $Y=910300
X1544 1557 1456 1550 1588 2 1 MXL2HS $T=690060 940920 1 0 $X=690060 $Y=935500
X1545 1558 1553 1582 1589 2 1 MXL2HS $T=690060 1021560 0 0 $X=690060 $Y=1021180
X1546 1546 1534 1580 1593 2 1 MXL2HS $T=690680 1051800 1 0 $X=690680 $Y=1046380
X1547 1569 1503 1516 1597 2 1 MXL2HS $T=692540 1011480 1 0 $X=692540 $Y=1006060
X1548 1595 1567 1579 1529 2 1 MXL2HS $T=699980 930840 0 180 $X=694400 $Y=925420
X1549 1605 1567 1596 1595 2 1 MXL2HS $T=700600 920760 1 180 $X=695020 $Y=920380
X1550 1607 1567 1574 1562 2 1 MXL2HS $T=701220 910680 1 180 $X=695640 $Y=910300
X1551 1573 1553 1600 1610 2 1 MXL2HS $T=695640 1031640 1 0 $X=695640 $Y=1026220
X1552 1589 1503 1584 1613 2 1 MXL2HS $T=696260 1001400 0 0 $X=696260 $Y=1001020
X1553 1577 1556 1592 1614 2 1 MXL2HS $T=696260 1051800 0 0 $X=696260 $Y=1051420
X1554 1532 129 1594 1615 2 1 MXL2HS $T=696260 1071960 1 0 $X=696260 $Y=1066540
X1555 1537 1602 1604 1618 2 1 MXL2HS $T=696880 951000 1 0 $X=696880 $Y=945580
X1556 1543 1553 1591 1619 2 1 MXL2HS $T=696880 1021560 0 0 $X=696880 $Y=1021180
X1557 1597 1503 1590 1632 2 1 MXL2HS $T=699360 1011480 1 0 $X=699360 $Y=1006060
X1558 1610 1553 1601 1634 2 1 MXL2HS $T=699980 1031640 0 0 $X=699980 $Y=1031260
X1559 1554 1621 1629 1637 2 1 MXL2HS $T=700600 981240 0 0 $X=700600 $Y=980860
X1560 1593 1556 1630 1641 2 1 MXL2HS $T=701840 1051800 1 0 $X=701840 $Y=1046380
X1561 1643 1567 1633 1607 2 1 MXL2HS $T=708040 910680 1 180 $X=702460 $Y=910300
X1562 1618 1602 1628 1645 2 1 MXL2HS $T=703700 951000 1 0 $X=703700 $Y=945580
X1563 1518 1635 1611 1651 2 1 MXL2HS $T=704320 961080 0 0 $X=704320 $Y=960700
X1564 1561 1635 1575 1653 2 1 MXL2HS $T=704940 971160 1 0 $X=704940 $Y=965740
X1565 1661 1567 1627 1605 2 1 MXL2HS $T=711760 930840 0 180 $X=706180 $Y=925420
X1566 1637 1621 1626 1667 2 1 MXL2HS $T=706800 981240 0 0 $X=706800 $Y=980860
X1567 1619 1649 1658 1669 2 1 MXL2HS $T=707420 1031640 1 0 $X=707420 $Y=1026220
X1568 1636 138 137 1587 2 1 MXL2HS $T=713620 900600 1 180 $X=708040 $Y=900220
X1569 1652 138 1656 1636 2 1 MXL2HS $T=714240 910680 0 180 $X=708660 $Y=905260
X1570 1614 1556 1668 1672 2 1 MXL2HS $T=708660 1051800 0 0 $X=708660 $Y=1051420
X1571 1613 1657 1671 1676 2 1 MXL2HS $T=709280 1001400 1 0 $X=709280 $Y=995980
X1572 1588 1602 1647 1679 2 1 MXL2HS $T=709900 940920 1 0 $X=709900 $Y=935500
X1573 1667 1635 1678 1686 2 1 MXL2HS $T=711140 971160 1 0 $X=711140 $Y=965740
X1574 1645 1602 1648 1689 2 1 MXL2HS $T=713000 951000 1 0 $X=713000 $Y=945580
X1575 1634 1649 1659 1690 2 1 MXL2HS $T=713000 1031640 0 0 $X=713000 $Y=1031260
X1576 1681 1657 1688 1696 2 1 MXL2HS $T=713620 991320 1 0 $X=713620 $Y=985900
X1577 1676 1657 1694 1681 2 1 MXL2HS $T=714240 991320 0 0 $X=714240 $Y=990940
X1578 1632 1649 1654 1697 2 1 MXL2HS $T=714240 1011480 0 0 $X=714240 $Y=1011100
X1579 1669 1649 1663 1698 2 1 MXL2HS $T=714240 1031640 1 0 $X=714240 $Y=1026220
X1580 1641 1556 1695 1701 2 1 MXL2HS $T=714860 1051800 0 0 $X=714860 $Y=1051420
X1581 1615 129 1665 1683 2 1 MXL2HS $T=715480 1071960 0 0 $X=715480 $Y=1071580
X1582 1704 1602 1692 1661 2 1 MXL2HS $T=721680 940920 0 180 $X=716100 $Y=935500
X1583 1686 1693 1699 1708 2 1 MXL2HS $T=716720 961080 0 0 $X=716720 $Y=960700
X1584 1696 1693 1718 1704 2 1 MXL2HS $T=720440 971160 1 0 $X=720440 $Y=965740
X1585 1697 1702 1719 1724 2 1 MXL2HS $T=721060 1011480 0 0 $X=721060 $Y=1011100
X1586 1708 145 1717 1652 2 1 MXL2HS $T=727260 920760 1 180 $X=721680 $Y=920380
X1587 140 1602 1713 1726 2 1 MXL2HS $T=721680 951000 1 0 $X=721680 $Y=945580
X1588 1651 1693 1710 1729 2 1 MXL2HS $T=722300 961080 0 0 $X=722300 $Y=960700
X1589 1683 129 1722 1730 2 1 MXL2HS $T=722300 1071960 0 0 $X=722300 $Y=1071580
X1590 1690 1649 1714 1733 2 1 MXL2HS $T=723540 1031640 1 0 $X=723540 $Y=1026220
X1591 1724 1702 1707 1737 2 1 MXL2HS $T=725400 1011480 1 0 $X=725400 $Y=1006060
X1592 1712 145 1741 1746 2 1 MXL2HS $T=727880 920760 0 0 $X=727880 $Y=920380
X1593 1746 145 1728 1643 2 1 MXL2HS $T=735940 920760 0 180 $X=730360 $Y=915340
X1594 1653 1693 1751 1760 2 1 MXL2HS $T=730360 971160 1 0 $X=730360 $Y=965740
X1595 1698 1649 1721 1763 2 1 MXL2HS $T=730360 1031640 1 0 $X=730360 $Y=1026220
X1596 148 145 1750 1765 2 1 MXL2HS $T=731600 910680 1 0 $X=731600 $Y=905260
X1597 1737 1322 1770 1776 2 1 MXL2HS $T=734700 1011480 0 0 $X=734700 $Y=1011100
X1598 150 145 152 1781 2 1 MXL2HS $T=735940 900600 0 0 $X=735940 $Y=900220
X1599 1689 1769 1779 1783 2 1 MXL2HS $T=736560 940920 1 0 $X=736560 $Y=935500
X1600 1701 1771 1715 1777 2 1 MXL2HS $T=736560 1051800 0 0 $X=736560 $Y=1051420
X1601 1730 1773 154 1784 2 1 MXL2HS $T=736560 1071960 0 0 $X=736560 $Y=1071580
X1602 1778 1782 1755 1774 2 1 MXL2HS $T=742760 1011480 0 180 $X=737180 $Y=1006060
X1603 1672 1771 1780 1786 2 1 MXL2HS $T=737180 1041720 0 0 $X=737180 $Y=1041340
X1604 1679 1769 1766 1791 2 1 MXL2HS $T=738420 930840 0 0 $X=738420 $Y=930460
X1605 1777 1773 1723 1793 2 1 MXL2HS $T=738420 1061880 0 0 $X=738420 $Y=1061500
X1606 1733 1782 1767 1778 2 1 MXL2HS $T=744620 1021560 0 180 $X=739040 $Y=1016140
X1607 1726 1769 1797 1804 2 1 MXL2HS $T=740900 951000 1 0 $X=740900 $Y=945580
X1608 1784 1773 159 1814 2 1 MXL2HS $T=743380 1071960 0 0 $X=743380 $Y=1071580
X1609 1791 1769 1794 1815 2 1 MXL2HS $T=744000 930840 0 0 $X=744000 $Y=930460
X1610 1760 1803 1809 1816 2 1 MXL2HS $T=744000 971160 1 0 $X=744000 $Y=965740
X1611 1786 1771 1812 1819 2 1 MXL2HS $T=744620 1041720 0 0 $X=744620 $Y=1041340
X1612 1763 1771 1799 1822 2 1 MXL2HS $T=745240 1041720 1 0 $X=745240 $Y=1036300
X1613 1793 1773 1789 1823 2 1 MXL2HS $T=745240 1061880 0 0 $X=745240 $Y=1061500
X1614 1781 1808 1817 1824 2 1 MXL2HS $T=745860 910680 0 0 $X=745860 $Y=910300
X1615 1776 1782 1818 1825 2 1 MXL2HS $T=745860 1021560 1 0 $X=745860 $Y=1016140
X1616 1729 1803 1788 1826 2 1 MXL2HS $T=746480 961080 0 0 $X=746480 $Y=960700
X1617 1774 1782 1795 1828 2 1 MXL2HS $T=746480 1001400 1 0 $X=746480 $Y=995980
X1618 1816 1803 1837 1842 2 1 MXL2HS $T=750820 971160 1 0 $X=750820 $Y=965740
X1619 1822 1771 1839 1846 2 1 MXL2HS $T=751440 1041720 1 0 $X=751440 $Y=1036300
X1620 1819 1771 1810 1847 2 1 MXL2HS $T=751440 1041720 0 0 $X=751440 $Y=1041340
X1621 1765 1808 1787 1848 2 1 MXL2HS $T=752060 930840 1 0 $X=752060 $Y=925420
X1622 1828 1782 1807 1849 2 1 MXL2HS $T=752060 1001400 1 0 $X=752060 $Y=995980
X1623 1826 1803 1820 1852 2 1 MXL2HS $T=752680 961080 0 0 $X=752680 $Y=960700
X1624 165 1773 167 1855 2 1 MXL2HS $T=753300 1071960 0 0 $X=753300 $Y=1071580
X1625 1824 1808 1829 1859 2 1 MXL2HS $T=755160 910680 0 0 $X=755160 $Y=910300
X1626 1847 1857 1836 1869 2 1 MXL2HS $T=757640 1031640 1 0 $X=757640 $Y=1026220
X1627 1860 1803 1838 168 2 1 MXL2HS $T=758880 971160 1 0 $X=758880 $Y=965740
X1628 1848 1769 1870 1880 2 1 MXL2HS $T=759500 940920 1 0 $X=759500 $Y=935500
X1629 1815 1864 1875 1882 2 1 MXL2HS $T=760120 930840 1 0 $X=760120 $Y=925420
X1630 1825 1857 1873 1883 2 1 MXL2HS $T=760120 1021560 1 0 $X=760120 $Y=1016140
X1631 1855 1865 1878 1885 2 1 MXL2HS $T=760120 1051800 0 0 $X=760120 $Y=1051420
X1632 1872 1871 1811 1860 2 1 MXL2HS $T=766320 981240 0 180 $X=760740 $Y=975820
X1633 1814 1773 169 1887 2 1 MXL2HS $T=760740 1071960 0 0 $X=760740 $Y=1071580
X1634 1889 1871 1861 1868 2 1 MXL2HS $T=766940 991320 1 180 $X=761360 $Y=990940
X1635 1846 1857 1881 1890 2 1 MXL2HS $T=761360 1041720 1 0 $X=761360 $Y=1036300
X1636 1868 1871 1858 1872 2 1 MXL2HS $T=768800 981240 1 180 $X=763220 $Y=980860
X1637 1880 1769 1898 1906 2 1 MXL2HS $T=765700 940920 1 0 $X=765700 $Y=935500
X1638 1823 1865 1892 1907 2 1 MXL2HS $T=765700 1061880 0 0 $X=765700 $Y=1061500
X1639 1852 1894 1905 1914 2 1 MXL2HS $T=766940 961080 1 0 $X=766940 $Y=955660
X1640 168 171 1910 172 2 1 MXL2HS $T=767560 900600 0 0 $X=767560 $Y=900220
X1641 1869 1899 1909 1919 2 1 MXL2HS $T=767560 1021560 0 0 $X=767560 $Y=1021180
X1642 1804 1894 1834 1922 2 1 MXL2HS $T=768180 951000 1 0 $X=768180 $Y=945580
X1643 1919 1899 1888 1889 2 1 MXL2HS $T=774380 1011480 0 180 $X=768800 $Y=1006060
X1644 1890 1913 1900 1931 2 1 MXL2HS $T=771900 1041720 1 0 $X=771900 $Y=1036300
X1645 1924 1864 1921 175 2 1 MXL2HS $T=772520 920760 1 0 $X=772520 $Y=915340
X1646 1932 1894 1902 1924 2 1 MXL2HS $T=778100 930840 0 180 $X=772520 $Y=925420
X1647 1842 1871 1929 1932 2 1 MXL2HS $T=772520 971160 1 0 $X=772520 $Y=965740
X1648 1936 171 1927 173 2 1 MXL2HS $T=778720 900600 1 180 $X=773140 $Y=900220
X1649 1849 1899 1891 1938 2 1 MXL2HS $T=773760 1001400 0 0 $X=773760 $Y=1001020
X1650 1883 1899 1935 1941 2 1 MXL2HS $T=774380 1021560 1 0 $X=774380 $Y=1016140
X1651 1922 1894 1911 1945 2 1 MXL2HS $T=775000 951000 1 0 $X=775000 $Y=945580
X1652 1882 1864 1926 177 2 1 MXL2HS $T=777480 920760 0 0 $X=777480 $Y=920380
X1653 1907 1944 1947 1957 2 1 MXL2HS $T=778100 1061880 0 0 $X=778100 $Y=1061500
X1654 1945 1950 1951 179 2 1 MXL2HS $T=779960 940920 1 0 $X=779960 $Y=935500
X1655 1938 1899 1960 1962 2 1 MXL2HS $T=779960 1001400 0 0 $X=779960 $Y=1001020
X1656 1954 1871 1930 1965 2 1 MXL2HS $T=781200 971160 0 0 $X=781200 $Y=970780
X1657 1941 1865 1939 1970 2 1 MXL2HS $T=781200 1021560 1 0 $X=781200 $Y=1016140
X1658 1885 1944 1895 1974 2 1 MXL2HS $T=781820 1051800 0 0 $X=781820 $Y=1051420
X1659 1887 1944 1948 1976 2 1 MXL2HS $T=783060 1071960 1 0 $X=783060 $Y=1066540
X1660 1977 182 1971 180 2 1 MXL2HS $T=789880 900600 1 180 $X=784300 $Y=900220
X1661 1965 1968 1956 183 2 1 MXL2HS $T=784300 920760 1 0 $X=784300 $Y=915340
X1662 1964 1980 1912 1972 2 1 MXL2HS $T=791120 991320 1 180 $X=785540 $Y=990940
X1663 1973 1899 1984 1964 2 1 MXL2HS $T=785540 1011480 1 0 $X=785540 $Y=1006060
X1664 1982 1950 1979 181 2 1 MXL2HS $T=791740 951000 1 180 $X=786160 $Y=950620
X1665 1991 1950 1978 1936 2 1 MXL2HS $T=792360 940920 0 180 $X=786780 $Y=935500
X1666 1972 1989 1916 1954 2 1 MXL2HS $T=792360 981240 1 180 $X=786780 $Y=980860
X1667 1962 1980 1917 1992 2 1 MXL2HS $T=786780 1001400 1 0 $X=786780 $Y=995980
X1668 1993 1865 1969 1973 2 1 MXL2HS $T=792360 1031640 1 180 $X=786780 $Y=1031260
X1669 1957 1944 1997 1993 2 1 MXL2HS $T=788640 1051800 0 0 $X=788640 $Y=1051420
X1670 1976 1944 1981 2008 2 1 MXL2HS $T=789880 1071960 1 0 $X=789880 $Y=1066540
X1671 2009 1989 1983 1982 2 1 MXL2HS $T=796080 971160 0 180 $X=790500 $Y=965740
X1672 1970 1865 2001 2011 2 1 MXL2HS $T=790500 1021560 1 0 $X=790500 $Y=1016140
X1673 1992 1989 1986 2016 2 1 MXL2HS $T=791740 991320 0 0 $X=791740 $Y=990940
X1674 1914 1950 1990 186 2 1 MXL2HS $T=792980 951000 0 0 $X=792980 $Y=950620
X1675 2016 1989 1996 2009 2 1 MXL2HS $T=799800 981240 1 180 $X=794220 $Y=980860
X1676 1931 1913 2002 2028 2 1 MXL2HS $T=794220 1041720 0 0 $X=794220 $Y=1041340
X1677 1859 1864 2030 187 2 1 MXL2HS $T=796080 910680 0 0 $X=796080 $Y=910300
X1678 2038 2034 2025 178 2 1 MXL2HS $T=802280 961080 1 180 $X=796700 $Y=960700
X1679 2039 2034 2022 2023 2 1 MXL2HS $T=802900 971160 0 180 $X=797320 $Y=965740
X1680 2041 2037 2004 2024 2 1 MXL2HS $T=802900 1031640 1 180 $X=797320 $Y=1031260
X1681 2008 2035 2042 2041 2 1 MXL2HS $T=799180 1051800 0 0 $X=799180 $Y=1051420
X1682 2052 1980 2026 2039 2 1 MXL2HS $T=806000 991320 1 180 $X=800420 $Y=990940
X1683 2023 1968 2020 188 2 1 MXL2HS $T=801040 920760 0 0 $X=801040 $Y=920380
X1684 2055 2034 2046 185 2 1 MXL2HS $T=807240 951000 1 180 $X=801660 $Y=950620
X1685 1974 2035 2056 2062 2 1 MXL2HS $T=802900 1051800 1 0 $X=802900 $Y=1046380
X1686 2053 1968 2063 192 2 1 MXL2HS $T=804760 930840 1 0 $X=804760 $Y=925420
X1687 2024 2054 2061 2071 2 1 MXL2HS $T=804760 1011480 0 0 $X=804760 $Y=1011100
X1688 2011 2054 2050 2072 2 1 MXL2HS $T=804760 1021560 1 0 $X=804760 $Y=1016140
X1689 2028 2035 2065 2073 2 1 MXL2HS $T=804760 1041720 1 0 $X=804760 $Y=1036300
X1690 1906 1968 2021 194 2 1 MXL2HS $T=814680 940920 0 180 $X=809100 $Y=935500
X1691 2073 2037 2080 2086 2 1 MXL2HS $T=809100 1031640 0 0 $X=809100 $Y=1031260
X1692 2071 1980 2079 2087 2 1 MXL2HS $T=809720 991320 1 0 $X=809720 $Y=985900
X1693 2086 2054 2076 2052 2 1 MXL2HS $T=815920 1011480 1 180 $X=810340 $Y=1011100
X1694 2062 2035 2077 2098 2 1 MXL2HS $T=813440 1041720 1 0 $X=813440 $Y=1036300
X1695 2091 2082 2094 197 2 1 MXL2HS $T=819640 951000 1 180 $X=814060 $Y=950620
X1696 2093 1968 2090 193 2 1 MXL2HS $T=820260 940920 0 180 $X=814680 $Y=935500
X1697 2104 2088 2074 2091 2 1 MXL2HS $T=820260 981240 1 180 $X=814680 $Y=980860
X1698 2087 2088 2100 2096 2 1 MXL2HS $T=815300 971160 1 0 $X=815300 $Y=965740
X1699 2106 1980 2112 2104 2 1 MXL2HS $T=819640 991320 0 0 $X=819640 $Y=990940
X1700 2072 2054 2108 2106 2 1 MXL2HS $T=825220 1011480 1 180 $X=819640 $Y=1011100
X1701 2098 2054 2097 2114 2 1 MXL2HS $T=819640 1021560 1 0 $X=819640 $Y=1016140
X1702 2096 2082 2111 196 2 1 MXL2HS $T=820260 951000 0 0 $X=820260 $Y=950620
X1703 2117 2088 2113 2038 2 1 MXL2HS $T=828320 971160 0 180 $X=822740 $Y=965740
X1704 2114 2054 2116 2122 2 1 MXL2HS $T=825840 1011480 0 0 $X=825840 $Y=1011100
X1705 2122 1980 2120 2117 2 1 MXL2HS $T=833280 991320 1 180 $X=827700 $Y=990940
X1706 2173 2171 229 2166 2 1 MXL2HS $T=873580 910680 0 180 $X=868000 $Y=905260
X1707 12 14 1 2 INV12CK $T=380060 1071960 0 0 $X=380060 $Y=1071580
X1708 12 20 1 2 INV12CK $T=388740 1051800 1 0 $X=388740 $Y=1046380
X1709 45 28 1 2 INV12CK $T=489800 900600 0 0 $X=489800 $Y=900220
X1710 795 340 1 2 INV12CK $T=504680 971160 0 0 $X=504680 $Y=970780
X1711 795 46 1 2 INV12CK $T=511500 961080 0 0 $X=511500 $Y=960700
X1712 795 49 1 2 INV12CK $T=525140 910680 0 0 $X=525140 $Y=910300
X1713 107 63 1 2 INV12CK $T=662780 971160 0 180 $X=652860 $Y=965740
X1714 107 1026 1 2 INV12CK $T=667740 951000 0 180 $X=657820 $Y=945580
X1715 1720 1583 1 2 INV12CK $T=724160 981240 0 0 $X=724160 $Y=980860
X1716 1720 102 1 2 INV12CK $T=731600 991320 0 0 $X=731600 $Y=990940
X1717 1720 147 1 2 INV12CK $T=745240 991320 0 0 $X=745240 $Y=990940
X1718 2314 2307 1 2 279 AN2 $T=967820 910680 1 0 $X=967820 $Y=905260
X1719 2134 2137 2132 1 2 ND2 $T=846300 910680 1 180 $X=844440 $Y=910300
X1720 220 2138 223 1 2 ND2 $T=848780 930840 0 0 $X=848780 $Y=930460
X1721 2155 2156 2143 1 2 ND2 $T=858700 930840 0 0 $X=858700 $Y=930460
X1722 230 2170 206 1 2 ND2 $T=871100 910680 1 180 $X=869240 $Y=910300
X1723 2174 2200 2148 1 2 ND2 $T=890320 930840 1 180 $X=888460 $Y=930460
X1724 2207 2209 214 1 2 ND2 $T=895280 940920 1 180 $X=893420 $Y=940540
X1725 2248 2262 2247 1 2 ND2 $T=920700 940920 0 0 $X=920700 $Y=940540
X1726 243 2280 265 1 2 ND2 $T=933100 900600 1 180 $X=931240 $Y=900220
X1727 2275 2287 2283 1 2 ND2 $T=938680 930840 1 180 $X=936820 $Y=930460
X1728 2303 275 2306 1 2 ND2 $T=957900 910680 1 0 $X=957900 $Y=905260
X1729 2305 2310 2297 1 2 ND2 $T=960380 930840 0 180 $X=958520 $Y=925420
X1730 2301 2307 2278 1 2 ND2 $T=961620 920760 0 180 $X=959760 $Y=915340
X1731 2296 2309 2297 1 2 ND2 $T=959760 930840 0 0 $X=959760 $Y=930460
X1732 2305 2312 2296 1 2 ND2 $T=964720 930840 1 180 $X=962860 $Y=930460
X1733 2313 276 2311 1 2 ND2 $T=967820 910680 1 180 $X=965960 $Y=910300
X1734 254 255 1 256 2 2249 OAI12HS $T=910160 900600 0 0 $X=910160 $Y=900220
X1735 2180 2248 1 2239 2 2253 OAI12HS $T=913880 940920 0 0 $X=913880 $Y=940540
X1736 2259 2252 1 2262 2 2269 OAI12HS $T=921940 951000 1 0 $X=921940 $Y=945580
X1737 2292 2294 1 2287 2 2297 OAI12HS $T=945500 940920 1 0 $X=945500 $Y=935500
X1738 273 276 1 2307 2 278 OAI12HS $T=965340 900600 0 0 $X=965340 $Y=900220
X1739 271 2303 1 2306 2 NR2T $T=956660 900600 0 0 $X=956660 $Y=900220
X1740 277 2313 1 2311 2 NR2T $T=968440 920760 0 180 $X=963480 $Y=915340
X1741 2150 1 2147 2151 2 2145 ND3 $T=857460 930840 0 180 $X=854980 $Y=925420
X1742 225 1 2134 2160 2 2136 ND3 $T=859940 910680 1 0 $X=859940 $Y=905260
X1743 2254 1 2251 2243 2 2257 ND3 $T=916980 961080 0 0 $X=916980 $Y=960700
X1744 2310 1 2309 2311 2 2312 ND3 $T=962240 930840 1 0 $X=962240 $Y=925420
X1745 2136 218 2140 2 1 XNR2HS $T=844440 900600 0 0 $X=844440 $Y=900220
X1746 2147 203 2142 2 1 XNR2HS $T=853120 930840 0 180 $X=847540 $Y=925420
X1747 210 2149 2135 2 1 XNR2HS $T=856840 920760 1 180 $X=851260 $Y=920380
X1748 206 2149 2132 2 1 XNR2HS $T=857460 910680 0 180 $X=851880 $Y=905260
X1749 222 212 2162 2 1 XNR2HS $T=861180 910680 0 0 $X=861180 $Y=910300
X1750 2149 214 2161 2 1 XNR2HS $T=869860 940920 0 180 $X=864280 $Y=935500
X1751 2165 2167 2171 2 1 XNR2HS $T=868000 920760 1 0 $X=868000 $Y=915340
X1752 235 2164 2180 2 1 XNR2HS $T=874820 940920 0 0 $X=874820 $Y=940540
X1753 2136 199 2183 2 1 XNR2HS $T=876680 910680 1 0 $X=876680 $Y=905260
X1754 222 2126 2188 2 1 XNR2HS $T=878540 920760 0 0 $X=878540 $Y=920380
X1755 215 2194 2193 2 1 XNR2HS $T=889080 910680 1 180 $X=883500 $Y=910300
X1756 2146 2194 2199 2 1 XNR2HS $T=889080 920760 1 0 $X=889080 $Y=915340
X1757 2141 2194 2212 2 1 XNR2HS $T=891560 930840 0 0 $X=891560 $Y=930460
X1758 2127 2207 2213 2 1 XNR2HS $T=891560 951000 1 0 $X=891560 $Y=945580
X1759 202 2194 2215 2 1 XNR2HS $T=900860 910680 1 180 $X=895280 $Y=910300
X1760 2222 2220 2216 2 1 XNR2HS $T=901480 951000 1 180 $X=895900 $Y=950620
X1761 2141 2207 2221 2 1 XNR2HS $T=896520 940920 0 0 $X=896520 $Y=940540
X1762 2126 2217 2223 2 1 XNR2HS $T=897760 930840 0 0 $X=897760 $Y=930460
X1763 202 245 2226 2 1 XNR2HS $T=899620 910680 1 0 $X=899620 $Y=905260
X1764 2152 2217 2232 2 1 XNR2HS $T=902100 940920 1 0 $X=902100 $Y=935500
X1765 2216 2225 2233 2 1 XNR2HS $T=902100 961080 0 0 $X=902100 $Y=960700
X1766 249 213 252 2 1 XNR2HS $T=905200 910680 1 0 $X=905200 $Y=905260
X1767 2233 2243 258 2 1 XNR2HS $T=909540 961080 0 0 $X=909540 $Y=960700
X1768 2239 2126 2265 2 1 XNR2HS $T=921320 930840 1 0 $X=921320 $Y=925420
X1769 2238 2208 2273 2 1 XNR2HS $T=926900 910680 0 0 $X=926900 $Y=910300
X1770 2269 2201 2277 2 1 XNR2HS $T=928760 951000 1 0 $X=928760 $Y=945580
X1771 2204 2264 2281 2 1 XNR2HS $T=931240 940920 1 0 $X=931240 $Y=935500
X1772 2273 2276 2282 2 1 XNR2HS $T=932480 910680 0 0 $X=932480 $Y=910300
X1773 2281 2275 2285 2 1 XNR2HS $T=936200 920760 0 0 $X=936200 $Y=920380
X1774 254 2170 2291 2 1 XNR2HS $T=939300 920760 1 0 $X=939300 $Y=915340
X1775 2291 2279 2293 2 1 XNR2HS $T=942400 920760 0 0 $X=942400 $Y=920380
X1776 2286 2277 2296 2 1 XNR2HS $T=943640 951000 1 0 $X=943640 $Y=945580
X1777 2289 2290 2304 2 1 XNR2HS $T=952940 951000 1 0 $X=952940 $Y=945580
X1778 2240 2304 2313 2 1 XNR2HS $T=961620 951000 1 0 $X=961620 $Y=945580
X1779 223 220 2134 1 2 XOR2H $T=852500 920760 1 0 $X=852500 $Y=915340
X1780 2305 2308 2303 1 2 XOR2H $T=962240 920760 1 180 $X=953560 $Y=920380
X1781 2296 2297 2308 1 2 XOR2H $T=955420 940920 1 0 $X=955420 $Y=935500
X1782 223 2 2145 220 1 NR2 $T=852500 930840 0 0 $X=852500 $Y=930460
X1783 2150 2 2155 2138 1 NR2 $T=857460 930840 1 180 $X=855600 $Y=930460
X1784 225 2 226 2153 1 NR2 $T=859940 900600 0 0 $X=859940 $Y=900220
X1785 218 2 2168 231 1 NR2 $T=868000 900600 0 0 $X=868000 $Y=900220
X1786 209 2 2172 2176 1 NR2 $T=873580 930840 0 0 $X=873580 $Y=930460
X1787 2167 2 2179 2165 1 NR2 $T=877300 920760 1 180 $X=875440 $Y=920380
X1788 231 2 2182 225 1 NR2 $T=880400 900600 1 180 $X=878540 $Y=900220
X1789 2175 2 2184 231 1 NR2 $T=879160 930840 1 0 $X=879160 $Y=925420
X1790 2150 2 2190 231 1 NR2 $T=882260 930840 1 0 $X=882260 $Y=925420
X1791 231 2 2189 2186 1 NR2 $T=884120 930840 1 180 $X=882260 $Y=930460
X1792 2188 2 2196 2144 1 NR2 $T=884740 920760 0 0 $X=884740 $Y=920380
X1793 2197 2 2202 2148 1 NR2 $T=889080 920760 1 180 $X=887220 $Y=920380
X1794 2208 2 2267 2238 1 NR2 $T=923800 920760 1 0 $X=923800 $Y=915340
X1795 243 2 2284 265 1 NR2 $T=938680 900600 0 0 $X=938680 $Y=900220
X1796 2289 2 2298 2290 1 NR2 $T=949220 940920 0 0 $X=949220 $Y=940540
X1797 2278 2 273 2301 1 NR2 $T=957280 920760 0 180 $X=955420 $Y=915340
X1798 2299 2 2288 1 274 NR2P $T=952940 910680 1 0 $X=952940 $Y=905260
X1799 2138 2143 1 2145 2144 2143 2 MOAI1 $T=847540 940920 1 0 $X=847540 $Y=935500
X1800 2193 2158 1 2163 239 2183 2 MOAI1 $T=887840 910680 0 180 $X=883500 $Y=905260
X1801 2158 2181 1 2174 2204 2206 2 MOAI1 $T=887840 940920 1 0 $X=887840 $Y=935500
X1802 2158 2203 1 2144 2208 2211 2 MOAI1 $T=890320 930840 1 0 $X=890320 $Y=925420
X1803 2158 2212 1 2174 2210 2197 2 MOAI1 $T=897760 920760 1 180 $X=893420 $Y=920380
X1804 2158 2199 1 2174 244 2218 2 MOAI1 $T=894660 920760 1 0 $X=894660 $Y=915340
X1805 236 2224 1 2219 2238 2226 2 MOAI1 $T=902720 920760 1 0 $X=902720 $Y=915340
X1806 2250 2241 1 2252 265 2260 2 MOAI1 $T=918840 910680 0 0 $X=918840 $Y=910300
X1807 2250 2270 1 2272 2279 2252 2 MOAI1 $T=927520 920760 0 0 $X=927520 $Y=920380
X1808 2290 2289 1 2302 2301 2298 2 MOAI1 $T=952320 940920 0 0 $X=952320 $Y=940540
X1809 2299 1 2288 272 2 ND2P $T=954180 900600 1 180 $X=950460 $Y=900220
X1810 2201 2286 2269 1 2 2290 MAO222 $T=938060 951000 1 0 $X=938060 $Y=945580
X1811 2170 2279 254 1 2 2300 MAO222 $T=946740 920760 1 0 $X=946740 $Y=915340
X1812 2240 2255 2 2209 2235 1 2263 FA1 $T=908300 951000 0 0 $X=908300 $Y=950620
X1813 260 2249 2 2182 2237 1 2276 FA1 $T=915120 900600 0 0 $X=915120 $Y=900220
X1814 268 2210 2 2266 266 1 2258 FA1 $T=935580 910680 0 180 $X=920080 $Y=905260
X1815 2275 2170 2 2184 2234 1 2286 FA1 $T=930620 930840 1 0 $X=930620 $Y=925420
X1816 270 2258 2 2293 2282 1 2299 FA1 $T=936820 910680 1 0 $X=936820 $Y=905260
X1817 2288 2285 2 2300 2274 1 2306 FA1 $T=942400 910680 0 0 $X=942400 $Y=910300
X1818 2305 2190 2 2295 2230 1 2289 FA1 $T=957900 930840 1 180 $X=942400 $Y=930460
X1819 2196 2202 2 1 243 OR2 $T=889700 920760 0 0 $X=889700 $Y=920380
X1820 2264 2204 2 1 2283 OR2 $T=939920 940920 0 180 $X=937440 $Y=935500
X1821 203 2172 2 2149 1 2169 AOI12HS $T=872960 930840 0 180 $X=868620 $Y=925420
X1822 2280 267 2 2284 1 269 AOI12HS $T=934340 900600 0 0 $X=934340 $Y=900220
X1823 209 206 211 2 1 XOR2HS $T=835760 910680 1 0 $X=835760 $Y=905260
X1824 220 206 224 2 1 XOR2HS $T=858700 900600 1 180 $X=853120 $Y=900220
X1825 209 210 232 2 1 XOR2HS $T=869240 920760 0 0 $X=869240 $Y=920380
X1826 2152 2194 2197 2 1 XOR2HS $T=884120 930840 1 0 $X=884120 $Y=925420
X1827 2181 2127 2203 2 1 XOR2HS $T=887840 940920 0 0 $X=887840 $Y=940540
X1828 213 2194 2205 2 1 XOR2HS $T=889080 910680 0 0 $X=889080 $Y=910300
X1829 213 245 247 2 1 XOR2HS $T=895900 900600 0 0 $X=895900 $Y=900220
X1830 2146 2217 2224 2 1 XOR2HS $T=898380 920760 0 0 $X=898380 $Y=920380
X1831 249 202 2241 2 1 XOR2HS $T=905200 910680 0 0 $X=905200 $Y=910300
X1832 2239 2127 2244 2 1 XOR2HS $T=907680 951000 1 0 $X=907680 $Y=945580
X1833 249 2146 2245 2 1 XOR2HS $T=908300 920760 0 0 $X=908300 $Y=920380
X1834 2242 2146 253 2 1 XOR2HS $T=914500 920760 0 180 $X=908920 $Y=915340
X1835 2127 2242 257 2 1 XOR2HS $T=908920 930840 0 0 $X=908920 $Y=930460
X1836 2141 2239 2247 2 1 XOR2HS $T=908920 940920 1 0 $X=908920 $Y=935500
X1837 2242 2126 261 2 1 XOR2HS $T=913880 920760 0 0 $X=913880 $Y=920380
X1838 2242 2141 263 2 1 XOR2HS $T=915120 930840 0 0 $X=915120 $Y=930460
X1839 2242 2152 264 2 1 XOR2HS $T=915740 930840 1 0 $X=915740 $Y=925420
X1840 2152 2239 2256 2 1 XOR2HS $T=921320 930840 0 0 $X=921320 $Y=930460
X1841 2253 2263 2268 2 1 XOR2HS $T=923180 961080 1 0 $X=923180 $Y=955660
X1842 2214 2268 2278 2 1 XOR2HS $T=930000 961080 1 0 $X=930000 $Y=955660
X1843 2138 2143 1 2145 2143 2154 2 MOAI1S $T=856220 940920 1 0 $X=856220 $Y=935500
X1844 236 2168 1 234 231 2166 2 MOAI1S $T=877920 900600 1 180 $X=874200 $Y=900220
X1845 2180 232 1 2169 2177 2167 2 MOAI1S $T=878540 930840 0 180 $X=874820 $Y=925420
X1846 2207 236 1 2219 2213 2220 2 MOAI1S $T=897760 951000 1 0 $X=897760 $Y=945580
X1847 2248 2244 1 2187 2252 2255 2 MOAI1S $T=913880 951000 1 0 $X=913880 $Y=945580
X1848 2208 2238 1 2271 2267 2274 2 MOAI1S $T=927520 920760 1 0 $X=927520 $Y=915340
X1849 2200 2201 2181 2 1 ND2S $T=889700 951000 0 180 $X=887840 $Y=945580
X1850 2207 2222 199 2 1 ND2S $T=900860 930840 1 0 $X=900860 $Y=925420
X1851 2214 2251 2253 2 1 ND2S $T=916360 961080 0 180 $X=914500 $Y=955660
X1852 2263 2254 2253 2 1 ND2S $T=917600 961080 1 0 $X=917600 $Y=955660
X1853 2214 2257 2263 2 1 ND2S $T=920700 961080 1 0 $X=920700 $Y=955660
X1854 204 205 1 2125 207 208 2 MOAI1H $T=830180 900600 0 0 $X=830180 $Y=900220
X1855 2134 2135 1 2139 219 2142 2 MOAI1H $T=843200 920760 1 0 $X=843200 $Y=915340
X1856 2165 2167 1 2173 237 2179 2 MOAI1H $T=873580 920760 1 0 $X=873580 $Y=915340
X1857 2215 2158 1 2205 242 2163 2 MOAI1H $T=896520 910680 0 180 $X=889080 $Y=905260
X1858 2248 2256 1 2261 2264 2252 2 MOAI1H $T=918220 940920 1 0 $X=918220 $Y=935500
X1859 2250 2245 1 2265 2266 2252 2 MOAI1H $T=920080 920760 0 0 $X=920080 $Y=920380
X1860 14 18 1 2 INV2 $T=380060 1071960 1 0 $X=380060 $Y=1066540
X1861 18 407 1 2 INV2 $T=405480 1041720 1 0 $X=405480 $Y=1036300
X1862 649 696 1 2 INV2 $T=479880 1011480 0 0 $X=479880 $Y=1011100
X1863 799 782 1 2 INV2 $T=505920 971160 0 180 $X=504060 $Y=965740
X1864 782 783 1 2 INV2 $T=507780 971160 1 0 $X=507780 $Y=965740
X1865 44 874 1 2 INV2 $T=527000 900600 0 0 $X=527000 $Y=900220
X1866 912 913 1 2 INV2 $T=536920 1041720 0 0 $X=536920 $Y=1041340
X1867 860 983 1 2 INV2 $T=551180 961080 0 0 $X=551180 $Y=960700
X1868 1156 1148 1 2 INV2 $T=592720 920760 1 180 $X=590860 $Y=920380
X1869 1156 1082 1 2 INV2 $T=591480 930840 1 0 $X=591480 $Y=925420
X1870 1170 1156 1 2 INV2 $T=595200 930840 0 0 $X=595200 $Y=930460
X1871 1108 1200 1 2 INV2 $T=598300 1051800 0 0 $X=598300 $Y=1051420
X1872 1200 1210 1 2 INV2 $T=602020 1051800 1 0 $X=602020 $Y=1046380
X1873 1200 76 1 2 INV2 $T=602020 1051800 0 0 $X=602020 $Y=1051420
X1874 144 1606 1 2 INV2 $T=724780 910680 1 0 $X=724780 $Y=905260
X1875 151 1762 1 2 INV2 $T=737800 981240 1 0 $X=737800 $Y=975820
X1876 158 1322 1 2 INV2 $T=742140 981240 1 180 $X=740280 $Y=980860
X1877 2134 2153 1 2 INV2 $T=856220 910680 0 0 $X=856220 $Y=910300
X1878 2157 2143 1 2 INV2 $T=859940 940920 1 180 $X=858080 $Y=940540
X1879 2161 2159 1 2 INV2 $T=864280 940920 0 180 $X=862420 $Y=935500
X1880 2164 2157 1 2 INV2 $T=865520 940920 1 180 $X=863660 $Y=940540
X1881 2157 2149 1 2 INV2 $T=869860 930840 0 0 $X=869860 $Y=930460
X1882 230 231 1 2 INV2 $T=870480 900600 0 0 $X=870480 $Y=900220
X1883 2164 2181 1 2 INV2 $T=878540 951000 1 0 $X=878540 $Y=945580
X1884 2192 205 1 2 INV2 $T=884120 900600 1 180 $X=882260 $Y=900220
X1885 2192 238 1 2 INV2 $T=884120 900600 0 0 $X=884120 $Y=900220
X1886 2180 259 1 2 INV2 $T=913260 910680 1 180 $X=911400 $Y=910300
X1887 254 2242 1 2 INV2 $T=915120 920760 1 0 $X=915120 $Y=915340
X1888 2192 2248 1 2 INV2 $T=915740 940920 1 0 $X=915740 $Y=935500
X1889 2192 2250 1 2 INV2 $T=918220 920760 1 0 $X=918220 $Y=915340
X1890 744 659 1 2 BUF2 $T=493520 971160 0 180 $X=490420 $Y=965740
X1891 783 768 1 2 BUF2 $T=517700 981240 0 0 $X=517700 $Y=980860
X1892 53 862 1 2 BUF2 $T=518940 1001400 0 0 $X=518940 $Y=1001020
X1893 819 787 1 2 BUF2 $T=527000 1061880 0 180 $X=523900 $Y=1056460
X1894 911 799 1 2 BUF2 $T=533200 971160 0 180 $X=530100 $Y=965740
X1895 871 792 1 2 BUF2 $T=533820 981240 0 180 $X=530720 $Y=975820
X1896 14 843 1 2 BUF2 $T=535060 1051800 1 0 $X=535060 $Y=1046380
X1897 843 894 1 2 BUF2 $T=536300 1011480 0 0 $X=536300 $Y=1011100
X1898 940 871 1 2 BUF2 $T=540640 991320 0 180 $X=537540 $Y=985900
X1899 787 943 1 2 BUF2 $T=540020 1071960 1 0 $X=540020 $Y=1066540
X1900 924 860 1 2 BUF2 $T=540640 951000 0 0 $X=540640 $Y=950620
X1901 931 917 1 2 BUF2 $T=549320 920760 1 180 $X=546220 $Y=920380
X1902 971 912 1 2 BUF2 $T=549320 1041720 1 180 $X=546220 $Y=1041340
X1903 894 955 1 2 BUF2 $T=548080 1021560 1 0 $X=548080 $Y=1016140
X1904 955 1012 1 2 BUF2 $T=557380 1021560 1 0 $X=557380 $Y=1016140
X1905 1007 971 1 2 BUF2 $T=567920 1031640 1 0 $X=567920 $Y=1026220
X1906 943 1108 1 2 BUF2 $T=573500 1061880 0 0 $X=573500 $Y=1061500
X1907 367 1069 1 2 BUF2 $T=579080 1061880 0 0 $X=579080 $Y=1061500
X1908 1076 1117 1 2 BUF2 $T=590860 940920 1 0 $X=590860 $Y=935500
X1909 1117 1207 1 2 BUF2 $T=600780 940920 1 0 $X=600780 $Y=935500
X1910 1117 1172 1 2 BUF2 $T=601400 951000 1 0 $X=601400 $Y=945580
X1911 1250 1170 1 2 BUF2 $T=619380 930840 1 180 $X=616280 $Y=930460
X1912 90 1250 1 2 BUF2 $T=629920 920760 1 180 $X=626820 $Y=920380
X1913 1305 1345 1 2 BUF2 $T=633640 930840 0 0 $X=633640 $Y=930460
X1914 1340 91 1 2 BUF2 $T=651620 1071960 0 180 $X=648520 $Y=1066540
X1915 1489 1439 1 2 BUF2 $T=672080 971160 0 180 $X=668980 $Y=965740
X1916 111 1438 1 2 BUF2 $T=675180 920760 0 180 $X=672080 $Y=915340
X1917 111 1507 1 2 BUF2 $T=674560 920760 0 0 $X=674560 $Y=920380
X1918 1434 1513 1 2 BUF2 $T=674560 1011480 1 0 $X=674560 $Y=1006060
X1919 1417 1463 1 2 BUF2 $T=675180 1051800 1 0 $X=675180 $Y=1046380
X1920 1417 121 1 2 BUF2 $T=676420 1061880 0 0 $X=676420 $Y=1061500
X1921 1581 1489 1 2 BUF2 $T=692540 961080 1 0 $X=692540 $Y=955660
X1922 1585 1666 1 2 BUF2 $T=710520 961080 0 0 $X=710520 $Y=960700
X1923 1606 139 1 2 BUF2 $T=715480 900600 0 0 $X=715480 $Y=900220
X1924 1625 1734 1 2 BUF2 $T=725400 1061880 1 0 $X=725400 $Y=1056460
X1925 1666 1736 1 2 BUF2 $T=730360 951000 0 0 $X=730360 $Y=950620
X1926 1734 1756 1 2 BUF2 $T=734700 1061880 1 0 $X=734700 $Y=1056460
X1927 1756 1840 1 2 BUF2 $T=758880 1051800 1 180 $X=755780 $Y=1051420
X1928 1840 1966 1 2 BUF2 $T=783680 1051800 1 0 $X=783680 $Y=1046380
X1929 1966 2033 1 2 BUF2 $T=798560 1041720 1 0 $X=798560 $Y=1036300
X1930 2153 2148 1 2 BUF2 $T=858080 910680 0 0 $X=858080 $Y=910300
X1931 248 2219 1 2 BUF2 $T=904580 910680 1 180 $X=901480 $Y=910300
X1932 259 2252 1 2 BUF2 $T=913880 910680 0 0 $X=913880 $Y=910300
X1933 262 2241 2180 2 2250 2246 1 AO22 $T=918840 910680 0 180 $X=913880 $Y=905260
X1934 18 367 1 2 INV3 $T=389980 1071960 0 0 $X=389980 $Y=1071580
X1935 20 43 1 2 INV3 $T=480500 1051800 1 0 $X=480500 $Y=1046380
X1936 782 744 1 2 INV3 $T=502820 971160 0 180 $X=500340 $Y=965740
X1937 913 819 1 2 INV3 $T=532580 1061880 0 180 $X=530100 $Y=1056460
X1938 983 911 1 2 INV3 $T=551180 971160 1 0 $X=551180 $Y=965740
X1939 1005 940 1 2 INV3 $T=556760 971160 1 180 $X=554280 $Y=970780
X1940 1027 1005 1 2 INV3 $T=560480 971160 1 180 $X=558000 $Y=970780
X1941 43 1585 1 2 INV3 $T=695640 991320 0 0 $X=695640 $Y=990940
X1942 222 2164 1 2 INV3 $T=866760 930840 0 0 $X=866760 $Y=930460
X1943 2239 2187 1 2 INV3 $T=909540 940920 0 0 $X=909540 $Y=940540
X1944 350 19 1 2 BUF6 $T=386880 1051800 0 0 $X=386880 $Y=1051420
X1945 1831 1867 1 2 BUF6 $T=763840 961080 0 0 $X=763840 $Y=960700
X1946 1867 1940 1 2 BUF6 $T=778100 961080 0 0 $X=778100 $Y=960700
X1947 1940 2003 1 2 BUF6 $T=796080 961080 1 180 $X=788640 $Y=960700
X1948 184 2012 1 2 BUF6 $T=797320 900600 0 0 $X=797320 $Y=900220
X1949 249 2239 1 2 BUF6 $T=907060 930840 1 0 $X=907060 $Y=925420
X1950 2148 1 2142 2133 221 2144 2 OAI22S $T=852500 910680 1 180 $X=848780 $Y=910300
X1951 2183 1 2153 2163 233 2162 2 OAI22S $T=877300 910680 1 180 $X=873580 $Y=910300
X1952 2188 1 2148 2144 240 2195 2 OAI22S $T=883500 920760 1 0 $X=883500 $Y=915340
X1953 2205 1 2153 2198 241 2163 2 OAI22S $T=892800 900600 1 180 $X=889080 $Y=900220
X1954 2213 1 2229 2219 2227 2221 2 OAI22S $T=906440 951000 0 180 $X=902720 $Y=945580
X1955 2223 1 2229 2219 2234 2231 2 OAI22S $T=903340 930840 1 0 $X=903340 $Y=925420
X1956 2221 1 2229 2219 2235 2232 2 OAI22S $T=903340 940920 0 0 $X=903340 $Y=940540
X1957 2232 1 2229 2219 2230 2223 2 OAI22S $T=907680 930840 1 180 $X=903960 $Y=930460
X1958 2226 1 251 248 2237 2228 2 OAI22S $T=908920 900600 1 180 $X=905200 $Y=900220
X1959 2225 2 2236 2189 2227 1 2214 FA1S $T=907680 961080 0 180 $X=895900 $Y=955660
X1960 18 343 1 2 INV4 $T=388120 1041720 1 0 $X=388120 $Y=1036300
X1961 14 22 1 2 INV4 $T=403000 1051800 0 0 $X=403000 $Y=1051420
X1962 20 44 1 2 INV4 $T=484840 1021560 0 0 $X=484840 $Y=1021180
X1963 2064 2101 1 2 INV4 $T=814060 1001400 0 0 $X=814060 $Y=1001020
X1964 2191 2192 1 2 INV4 $T=884740 940920 1 0 $X=884740 $Y=935500
X1965 2185 2187 2181 235 1 2 NR3HP $T=880400 940920 0 0 $X=880400 $Y=940540
X1966 1762 149 1 153 2 OR2T $T=734080 981240 0 0 $X=734080 $Y=980860
X1967 1796 151 1 155 2 OR2T $T=747100 981240 0 180 $X=740900 $Y=975820
X1968 2178 2185 1 2191 2 OR2T $T=878540 940920 1 0 $X=878540 $Y=935500
X1969 209 2177 2175 2176 2 2181 1 AOI13HS $T=876680 930840 0 0 $X=876680 $Y=930460
X1970 209 2 2176 2164 2178 1 NR3 $T=876060 940920 0 180 $X=872960 $Y=935500
X1971 2140 2139 2137 1 2 217 OA12 $T=850020 910680 0 180 $X=846300 $Y=905260
X1972 2149 2163 2160 1 2 228 OA12 $T=868000 910680 0 180 $X=864280 $Y=905260
X1973 2159 2139 1 2162 2165 2148 2 OAI22H $T=861800 920760 0 0 $X=861800 $Y=920380
X1974 2148 2159 1 2151 227 2156 2 OAI112H $T=865520 930840 0 180 $X=858080 $Y=925420
X1975 1994 1583 2129 2146 1 2 QDFFRBP $T=838860 920760 0 0 $X=838860 $Y=920380
X1976 1995 1583 2121 2 1 214 QDFFRBS $T=828320 930840 0 0 $X=828320 $Y=930460
X1977 1606 1529 1 96 134 2 1562 132 136 OAI222S $T=699360 910680 1 0 $X=699360 $Y=905260
X1978 1606 1605 1 1636 134 2 1643 142 136 OAI222S $T=714240 910680 1 0 $X=714240 $Y=905260
X1979 1606 1704 1 1708 134 2 1712 1711 136 OAI222S $T=726640 920760 0 180 $X=721060 $Y=915340
X1980 1963 1965 1 1882 1915 2 1977 1994 1988 OAI222S $T=784300 920760 0 0 $X=784300 $Y=920380
X1981 1963 181 1 1924 1915 2 1936 1995 1988 OAI222S $T=785540 930840 1 0 $X=785540 $Y=925420
X1982 2007 183 1 177 2000 2 180 2006 184 OAI222S $T=796080 900600 1 180 $X=790500 $Y=900220
X1983 1963 1982 1 1932 2013 2 1991 2049 1988 OAI222S $T=792980 940920 0 0 $X=792980 $Y=940540
X1984 2007 178 1 179 1915 2 185 2032 2012 OAI222S $T=793600 920760 1 0 $X=793600 $Y=915340
X1985 2007 188 1 187 2000 2 189 2058 2012 OAI222S $T=800420 910680 1 0 $X=800420 $Y=905260
X1986 2007 2023 1 1859 2000 2 190 2060 2012 OAI222S $T=801040 920760 1 0 $X=801040 $Y=915340
X1987 1963 2038 1 1945 2013 2 2055 2067 1988 OAI222S $T=810960 951000 0 180 $X=805380 $Y=945580
X1988 2007 196 1 186 2000 2 192 2066 2012 OAI222S $T=812820 920760 1 180 $X=807240 $Y=920380
X1989 2007 197 1 194 2000 2 193 2075 2012 OAI222S $T=813440 920760 0 180 $X=807860 $Y=915340
X1990 1963 2096 1 1914 2013 2 2053 2084 1988 OAI222S $T=818400 951000 0 180 $X=812820 $Y=945580
X1991 1963 2091 1 1906 2013 2 2093 2099 1988 OAI222S $T=820260 940920 1 180 $X=814680 $Y=940540
X1992 473 28 453 2 1 514 518 28 525 551 293 ICV_12 $T=425940 940920 0 0 $X=425940 $Y=940540
X1993 497 28 343 2 1 531 490 28 460 577 293 ICV_12 $T=430900 971160 0 0 $X=430900 $Y=970780
X1994 613 340 643 2 1 647 657 340 643 677 293 ICV_12 $T=460660 1041720 0 0 $X=460660 $Y=1041340
X1995 662 340 42 2 1 706 712 340 42 760 293 ICV_12 $T=473060 1071960 0 0 $X=473060 $Y=1071580
X1996 769 340 746 2 1 811 818 46 746 844 293 ICV_12 $T=497240 1021560 1 0 $X=497240 $Y=1016140
X1997 48 49 47 2 1 55 57 49 856 58 293 ICV_12 $T=502820 900600 0 0 $X=502820 $Y=900220
X1998 822 46 750 2 1 857 863 46 843 886 293 ICV_12 $T=509640 1041720 1 0 $X=509640 $Y=1036300
X1999 823 46 42 2 1 859 864 46 891 906 293 ICV_12 $T=509640 1071960 0 0 $X=509640 $Y=1071580
X2000 830 46 871 2 1 848 899 46 871 925 293 ICV_12 $T=518940 991320 0 0 $X=518940 $Y=990940
X2001 920 46 891 2 1 960 968 63 891 1020 293 ICV_12 $T=536300 1071960 0 0 $X=536300 $Y=1071580
X2002 1019 46 1027 2 1 1065 1071 63 1027 1126 293 ICV_12 $T=558620 981240 1 0 $X=558620 $Y=975820
X2003 1025 63 891 2 1 1070 1078 63 367 1112 293 ICV_12 $T=559860 1071960 0 0 $X=559860 $Y=1071580
X2004 1174 1026 1207 2 1 1223 1225 1026 1207 1267 293 ICV_12 $T=595200 930840 1 0 $X=595200 $Y=925420
X2005 1169 74 1207 2 1 1224 1239 74 1259 1265 293 ICV_12 $T=597060 910680 0 0 $X=597060 $Y=910300
X2006 1184 63 1217 2 1 1234 1241 1026 1217 1276 293 ICV_12 $T=597060 981240 1 0 $X=597060 $Y=975820
X2007 1266 1026 1321 2 1 1309 1334 1026 1321 1380 293 ICV_12 $T=621860 971160 1 0 $X=621860 $Y=965740
X2008 1315 63 1344 2 1 1343 1360 63 1344 1410 293 ICV_12 $T=628060 1021560 0 0 $X=628060 $Y=1021180
X2009 1402 1026 1438 2 1 1430 1448 1026 1438 1483 293 ICV_12 $T=650380 930840 0 0 $X=650380 $Y=930460
X2010 1409 1026 1439 2 1 1443 1450 102 1439 1478 293 ICV_12 $T=650380 981240 1 0 $X=650380 $Y=975820
X2011 1395 1026 1439 2 1 1453 1460 102 1439 1502 293 ICV_12 $T=651620 971160 0 0 $X=651620 $Y=970780
X2012 1408 1026 1439 2 1 1452 1465 1026 1439 1504 293 ICV_12 $T=652240 961080 0 0 $X=652240 $Y=960700
X2013 1579 1583 1603 2 1 1608 1627 1583 1603 1677 293 ICV_12 $T=690680 930840 0 0 $X=690680 $Y=930460
X2014 1548 1026 1581 2 1 1572 1626 102 1585 1675 293 ICV_12 $T=690680 981240 1 0 $X=690680 $Y=975820
X2015 1659 102 1624 2 1 1709 1714 102 1734 1748 293 ICV_12 $T=709900 1041720 1 0 $X=709900 $Y=1036300
X2016 1721 102 1744 2 1 1764 1767 102 1744 1798 293 ICV_12 $T=724160 1021560 0 0 $X=724160 $Y=1021180
X2017 1861 147 1893 2 1 1901 1917 147 1893 1959 293 ICV_12 $T=759500 1001400 1 0 $X=759500 $Y=995980
X2018 1898 1583 1933 2 1 1928 1951 1583 1933 1999 293 ICV_12 $T=768800 940920 0 0 $X=768800 $Y=940540
X2019 1927 127 19 2 1 1952 1971 127 19 1998 293 ICV_12 $T=774380 910680 1 0 $X=774380 $Y=905260
X2020 191 127 195 2 1 198 2006 127 200 203 293 ICV_12 $T=806620 900600 0 0 $X=806620 $Y=900220
X2021 917 2 1 64 BUF3 $T=548700 900600 0 0 $X=548700 $Y=900220
X2022 1012 2 1 1027 BUF3 $T=568540 991320 0 0 $X=568540 $Y=990940
X2023 1045 2 1 1076 BUF3 $T=584040 920760 1 0 $X=584040 $Y=915340
X2024 1736 2 1 1831 BUF3 $T=748340 951000 0 0 $X=748340 $Y=950620
X2025 2003 2 1 2019 BUF3 $T=805380 991320 1 0 $X=805380 $Y=985900
X2026 2019 2064 1 2 INV6 $T=809100 1001400 1 180 $X=804140 $Y=1001020
X2027 388 6 372 2 1 419 419 436 293 ICV_13 $T=399900 981240 0 0 $X=399900 $Y=980860
X2028 424 6 453 2 1 462 462 438 293 ICV_13 $T=411680 940920 0 0 $X=411680 $Y=940540
X2029 435 6 453 2 1 493 493 446 293 ICV_13 $T=419120 971160 1 0 $X=419120 $Y=965740
X2030 494 28 470 2 1 532 532 543 293 ICV_13 $T=430280 920760 0 0 $X=430280 $Y=920380
X2031 500 340 523 2 1 535 535 554 293 ICV_13 $T=431520 1001400 0 0 $X=431520 $Y=1001020
X2032 476 340 520 2 1 536 536 485 293 ICV_13 $T=431520 1041720 0 0 $X=431520 $Y=1041340
X2033 603 28 563 2 1 670 670 572 293 ICV_13 $T=463140 961080 0 0 $X=463140 $Y=960700
X2034 851 49 874 2 1 892 892 904 293 ICV_13 $T=518320 930840 1 0 $X=518320 $Y=925420
X2035 993 46 1012 2 1 1041 1041 1031 293 ICV_13 $T=553660 1011480 1 0 $X=553660 $Y=1006060
X2036 1216 1026 1172 2 1 1260 1260 1242 293 ICV_13 $T=604500 951000 0 0 $X=604500 $Y=950620
X2037 1379 63 1384 2 1 1426 1426 1335 293 ICV_13 $T=644180 1041720 1 0 $X=644180 $Y=1036300
X2038 1549 1026 1581 2 1 1623 1623 1562 293 ICV_13 $T=690680 971160 0 0 $X=690680 $Y=970780
X2039 1596 1026 1603 2 1 1682 1682 1605 293 ICV_13 $T=703080 920760 0 0 $X=703080 $Y=920380
X2040 1654 102 1624 2 1 1706 1706 1632 293 ICV_13 $T=709280 1011480 1 0 $X=709280 $Y=1006060
X2041 1895 147 1923 2 1 1942 1942 1885 293 ICV_13 $T=767560 1051800 0 0 $X=767560 $Y=1051420
X2042 1912 147 1893 2 1 1955 1955 1964 293 ICV_13 $T=770660 991320 0 0 $X=770660 $Y=990940
X2043 2026 147 2019 2 1 2070 2057 2071 293 ICV_13 $T=797940 1001400 1 0 $X=797940 $Y=995980
X2044 2025 1583 2078 2 1 2089 2089 2038 293 ICV_13 $T=803520 961080 0 0 $X=803520 $Y=960700
X2045 333 340 361 2 1 369 374 340 361 406 293 ICV_14 $T=382540 1011480 1 0 $X=382540 $Y=1006060
X2046 495 340 520 2 1 528 540 340 520 567 293 ICV_14 $T=430280 1061880 0 0 $X=430280 $Y=1061500
X2047 511 340 460 2 1 555 559 340 585 596 293 ICV_14 $T=435860 991320 1 0 $X=435860 $Y=985900
X2048 660 340 696 2 1 703 709 340 746 759 293 ICV_14 $T=472440 1021560 1 0 $X=472440 $Y=1016140
X2049 679 340 694 2 1 720 727 340 733 757 293 ICV_14 $T=475540 1001400 0 0 $X=475540 $Y=1001020
X2050 710 340 750 2 1 762 756 340 750 815 293 ICV_14 $T=485460 1041720 0 0 $X=485460 $Y=1041340
X2051 813 46 750 2 1 850 861 46 843 902 293 ICV_14 $T=508400 1051800 1 0 $X=508400 $Y=1046380
X2052 820 46 843 2 1 858 866 46 894 872 293 ICV_14 $T=509640 1011480 0 0 $X=509640 $Y=1011100
X2053 910 46 939 2 1 954 961 46 939 1004 293 ICV_14 $T=533200 961080 1 0 $X=533200 $Y=955660
X2054 936 49 931 2 1 982 989 49 931 1034 293 ICV_14 $T=540020 930840 1 0 $X=540020 $Y=925420
X2055 947 46 940 2 1 988 995 46 1012 1053 293 ICV_14 $T=542500 991320 0 0 $X=542500 $Y=990940
X2056 1000 46 1013 2 1 1049 1058 46 1013 1094 293 ICV_14 $T=555520 1051800 1 0 $X=555520 $Y=1046380
X2057 1043 49 1076 2 1 1096 1103 1026 1076 1146 293 ICV_14 $T=565440 930840 1 0 $X=565440 $Y=925420
X2058 1122 63 1149 2 1 1163 1167 63 1149 1218 293 ICV_14 $T=581560 991320 0 0 $X=581560 $Y=990940
X2059 1123 63 367 2 1 1159 73 63 1213 79 293 ICV_14 $T=583420 1071960 0 0 $X=583420 $Y=1071580
X2060 1303 1026 1321 2 1 1346 1355 1026 1321 1400 293 ICV_14 $T=625580 951000 0 0 $X=625580 $Y=950620
X2061 1580 102 130 2 1 1612 1630 102 130 1664 293 ICV_14 $T=690680 1041720 0 0 $X=690680 $Y=1041340
X2062 2001 147 2033 2 1 2045 2050 147 2033 2092 293 ICV_14 $T=791740 1021560 0 0 $X=791740 $Y=1021180
X2063 2022 1583 2003 2 1 2069 2074 1583 2003 2107 293 ICV_14 $T=797320 981240 1 0 $X=797320 $Y=975820
X2064 2012 1 1988 2 BUF4CK $T=794840 920760 0 0 $X=794840 $Y=920380
X2065 1 2 496 468 512 475 504 439 293 ICV_15 $T=431520 1031640 0 180 $X=430280 $Y=1026220
X2066 1 2 705 695 732 659 697 695 293 ICV_15 $T=484220 981240 1 180 $X=482980 $Y=980860
X2067 1 2 811 801 832 797 818 802 293 ICV_15 $T=509020 1021560 1 180 $X=507780 $Y=1021180
X2068 1 2 827 805 836 768 830 805 293 ICV_15 $T=510880 991320 1 180 $X=509640 $Y=990940
X2069 1 2 844 832 868 797 855 832 293 ICV_15 $T=517700 1021560 1 180 $X=516460 $Y=1021180
X2070 1 2 880 868 901 900 889 868 293 ICV_15 $T=527000 1021560 1 180 $X=525760 $Y=1021180
X2071 1 2 942 915 965 924 935 915 293 ICV_15 $T=541880 951000 0 180 $X=540640 $Y=945580
X2072 1 2 960 930 981 943 968 930 293 ICV_15 $T=545600 1071960 0 180 $X=544360 $Y=1066540
X2073 1 2 976 965 987 924 963 965 293 ICV_15 $T=549940 951000 0 180 $X=548700 $Y=945580
X2074 1 2 988 969 1011 862 995 969 293 ICV_15 $T=552420 1001400 0 180 $X=551180 $Y=995980
X2075 1 2 1004 977 1029 992 1017 977 293 ICV_15 $T=556140 961080 1 180 $X=554900 $Y=960700
X2076 1 2 1049 1032 1073 971 1058 999 293 ICV_15 $T=566060 1041720 1 180 $X=564820 $Y=1041340
X2077 1 2 1065 1046 1089 1042 1071 1046 293 ICV_15 $T=569780 971160 1 180 $X=568540 $Y=970780
X2078 1 2 1070 1035 1093 943 1078 1052 293 ICV_15 $T=570400 1071960 0 180 $X=569160 $Y=1066540
X2079 1 2 1313 1301 1332 1298 1320 1301 293 ICV_15 $T=628680 971160 1 180 $X=627440 $Y=970780
X2080 1 2 1443 1411 1467 1403 1450 1444 293 ICV_15 $T=659680 981240 1 180 $X=658440 $Y=980860
X2081 1 2 1830 1791 1783 1808 1805 162 293 ICV_15 $T=751440 930840 1 180 $X=750200 $Y=930460
X2082 56 795 1 2 INV8CK $T=514600 910680 0 0 $X=514600 $Y=910300
X2083 143 1720 1 2 INV8CK $T=723540 971160 0 0 $X=723540 $Y=970780
X2084 64 1045 1 2 BUF4 $T=564820 900600 0 0 $X=564820 $Y=900220
X2085 12 16 1 2 INV4CK $T=381300 1051800 0 0 $X=381300 $Y=1051420
.ENDS
***************************************
.SUBCKT XOR3 I2 I1 I3 VCC GND O
** N=7 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ND3P I1 O I2 I3 GND VCC
** N=7 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OR2P I2 I1 O GND VCC
** N=6 EP=5 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT NR2F I1 VCC GND I2 O
** N=6 EP=5 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT DFFRBP D CK RB Q QB GND VCC
** N=8 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT INV3CK I GND VCC O
** N=5 EP=4 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT INV12 O I GND VCC
** N=5 EP=4 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OAI12HP B2 B1 GND A1 O VCC
** N=7 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OAI112HS C2 C1 GND B1 O A1 VCC
** N=8 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT DFFRBN D CK RB Q GND VCC QB
** N=8 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ND3HT I3 GND I2 I1 VCC O
** N=7 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AOI22S A1 B1 O B2 GND A2 VCC
** N=8 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT NR3H O I3 I2 I1 VCC GND
** N=7 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT BUF1CK I GND VCC O
** N=5 EP=4 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT BUF8CK I GND VCC O
** N=5 EP=4 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OAI12H B2 B1 GND A1 O VCC
** N=7 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ND3S I3 GND I2 O I1 VCC
** N=7 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AOI12H B2 B1 VCC O A1 GND
** N=7 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT HA1 A B C GND VCC S
** N=7 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_17 1 2 3 4 5 6 7 8 9
** N=9 EP=9 IP=12 FDC=0
X0 1 2 3 4 5 6 QDFFRBN $T=0 0 0 0 $X=0 $Y=-380
X1 7 4 8 5 INV1S $T=11780 0 0 0 $X=11780 $Y=-380
.ENDS
***************************************
.SUBCKT ICV_18 1 2 3 4 5 6 7 8 9 10 11
** N=11 EP=11 IP=14 FDC=0
X0 1 2 3 4 5 6 MXL2HS $T=-5580 0 0 0 $X=-5580 $Y=-380
X1 7 8 9 10 5 6 MXL2HS $T=0 0 0 0 $X=0 $Y=-380
.ENDS
***************************************
.SUBCKT ND2T I2 GND I1 O VCC
** N=6 EP=5 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT XNR3 I2 I1 I3 VCC GND O
** N=7 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MXL2H B S OB A GND VCC
** N=7 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT BUF6CK I GND O VCC
** N=5 EP=4 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT INV6CK I O GND VCC
** N=5 EP=4 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AOI22H A2 A1 VCC B1 O B2 GND
** N=8 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MAOI1H B1 B2 A2 A1 VCC GND O
** N=8 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MXL2HP B S OB A GND VCC
** N=7 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT BUF3CK I GND VCC O
** N=5 EP=4 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT XNR2H I2 O I1 GND VCC
** N=6 EP=5 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OA12P B2 B1 A1 O GND VCC
** N=7 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OAI12HT B2 B1 GND A1 O VCC
** N=7 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT DFFRBS D CK RB Q GND VCC QB
** N=8 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_19 1 2 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21
+ 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41
+ 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61
+ 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81
+ 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101
+ 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121
+ 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140 141
+ 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161
+ 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180 181
+ 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200 201
+ 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220 221
+ 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240 241
+ 242 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 259 260 261
+ 262 263 264 265 266 267 268 269 270 271 272 273 274 275 276 277 278 279 280 281
+ 282 283 284 285 286 287 288 289 290 291 292 293 294 295 296 297 298 299 300 301
+ 302 303 304 305 306 307 308 309 310 311 312 313 314 315 316 317 318 319 320 321
+ 322 323 324 325 326 327 328 329 330 331 332 333 334 335 336 337 338 339 340 341
+ 342 343 344 345 346 347 348 349 350 351 352 353 354 355 356 357 358 359 360 361
+ 362 363 364 365 366 367 368 369 370 371 372 373 374 375 376 377 378 379 380 381
+ 382 383 384 385 386 387 388 389 390 391 392 393 394 395 396 397 398 399 400 401
+ 402 403 404 405 406 407 408 409 410 411 412 413 414 415 416 417 418 419 420 421
+ 422 423 424 425 426 427 428 429 430 431 432 433 434 435 436 437 438 439 440 441
+ 442 443 444 445 446 447 448 449 450 451 452 453 454 455 456 457 458 459 460 461
+ 462 463 464 465 466 467 468 469 470 471 472 473 474 475 476 477 478 479 480 481
+ 482 483 484 485 486 487 488 489 490 491 492 493 494 495 496 497 498 499 500 501
+ 502 503 504 505 506 507 508 509 510 511 512 513 514 515 516 517 518 519 520 521
+ 522 523 524 525 526 527 528 529 530 531 532 533 534 535 536 537 538 539 540 541
+ 542 543 544 545 546 547 548 549 550 551 552 553 554 555 556 557 558 559 560 561
+ 562 563 564 565 566 567 568 569 570 571 572 589
** N=3753 EP=572 IP=21188 FDC=0
X0 1049 1 2 75 BUF1S $T=425320 729240 0 0 $X=425320 $Y=728860
X1 2437 1 2 2397 BUF1S $T=745860 819960 1 0 $X=745860 $Y=814540
X2 2408 1 2 2441 BUF1S $T=747100 749400 1 0 $X=747100 $Y=743980
X3 3350 1 2 3479 BUF1S $T=936820 769560 1 0 $X=936820 $Y=764140
X4 572 1 2 571 BUF1S $T=1129640 789720 0 180 $X=1127160 $Y=784300
X5 32 2 1 756 BUF1 $T=370760 900600 1 0 $X=370760 $Y=895180
X6 42 2 1 28 BUF1 $T=386260 900600 0 180 $X=383780 $Y=895180
X7 886 2 1 894 BUF1 $T=391220 850200 0 180 $X=388740 $Y=844780
X8 858 2 1 42 BUF1 $T=388740 880440 1 0 $X=388740 $Y=875020
X9 824 2 1 935 BUF1 $T=393700 870360 0 0 $X=393700 $Y=869980
X10 883 2 1 914 BUF1 $T=399280 850200 1 0 $X=399280 $Y=844780
X11 858 2 1 883 BUF1 $T=401760 860280 1 180 $X=399280 $Y=859900
X12 960 2 1 878 BUF1 $T=404860 739320 0 180 $X=402380 $Y=733900
X13 883 2 1 971 BUF1 $T=403000 860280 0 0 $X=403000 $Y=859900
X14 886 2 1 992 BUF1 $T=406720 850200 1 0 $X=406720 $Y=844780
X15 992 2 1 943 BUF1 $T=409820 840120 1 180 $X=407340 $Y=839740
X16 56 2 1 1017 BUF1 $T=411060 729240 1 0 $X=411060 $Y=723820
X17 64 2 1 858 BUF1 $T=414780 880440 0 180 $X=412300 $Y=875020
X18 1048 2 1 984 BUF1 $T=425940 819960 1 180 $X=423460 $Y=819580
X19 1110 2 1 1074 BUF1 $T=438340 809880 1 180 $X=435860 $Y=809500
X20 1029 2 1 1133 BUF1 $T=439580 809880 0 0 $X=439580 $Y=809500
X21 1130 2 1 76 BUF1 $T=443300 890520 0 180 $X=440820 $Y=885100
X22 1090 2 1 1097 BUF1 $T=448260 850200 0 180 $X=445780 $Y=844780
X23 1130 2 1 1129 BUF1 $T=446400 880440 0 0 $X=446400 $Y=880060
X24 1097 2 1 1122 BUF1 $T=447640 860280 1 0 $X=447640 $Y=854860
X25 1090 2 1 1163 BUF1 $T=448260 840120 0 0 $X=448260 $Y=839740
X26 1130 2 1 97 BUF1 $T=448880 890520 1 0 $X=448880 $Y=885100
X27 1172 2 1 1110 BUF1 $T=453840 799800 1 180 $X=451360 $Y=799420
X28 1126 2 1 1197 BUF1 $T=461280 830040 1 0 $X=461280 $Y=824620
X29 113 2 1 1220 BUF1 $T=468720 809880 1 0 $X=468720 $Y=804460
X30 1241 2 1 1262 BUF1 $T=474920 779640 0 0 $X=474920 $Y=779260
X31 1238 2 1 1287 BUF1 $T=478020 850200 0 0 $X=478020 $Y=849820
X32 1282 2 1 1241 BUF1 $T=481120 779640 1 180 $X=478640 $Y=779260
X33 1226 2 1 1299 BUF1 $T=485460 870360 1 0 $X=485460 $Y=864940
X34 1308 2 1 1227 BUF1 $T=488560 809880 1 180 $X=486080 $Y=809500
X35 1250 2 1 1337 BUF1 $T=488560 840120 0 0 $X=488560 $Y=839740
X36 1220 2 1 1367 BUF1 $T=496620 749400 0 0 $X=496620 $Y=749020
X37 1337 2 1 1368 BUF1 $T=503440 840120 1 180 $X=500960 $Y=839740
X38 1337 2 1 1395 BUF1 $T=502820 840120 1 0 $X=502820 $Y=834700
X39 1396 2 1 1251 BUF1 $T=506540 759480 0 180 $X=504060 $Y=754060
X40 1337 2 1 1308 BUF1 $T=506540 830040 0 180 $X=504060 $Y=824620
X41 146 2 1 1346 BUF1 $T=510260 729240 1 180 $X=507780 $Y=728860
X42 1367 2 1 1286 BUF1 $T=509020 749400 0 0 $X=509020 $Y=749020
X43 1414 2 1 1360 BUF1 $T=512120 789720 1 180 $X=509640 $Y=789340
X44 1422 2 1 1315 BUF1 $T=513360 880440 0 180 $X=510880 $Y=875020
X45 1419 2 1 1396 BUF1 $T=514600 759480 1 0 $X=514600 $Y=754060
X46 1396 2 1 1444 BUF1 $T=515840 769560 0 0 $X=515840 $Y=769180
X47 1382 2 1 1325 BUF1 $T=516460 749400 1 0 $X=516460 $Y=743980
X48 1414 2 1 1458 BUF1 $T=518320 799800 0 0 $X=518320 $Y=799420
X49 1395 2 1 1414 BUF1 $T=518320 819960 1 0 $X=518320 $Y=814540
X50 146 2 1 1419 BUF1 $T=520800 739320 0 0 $X=520800 $Y=738940
X51 1419 2 1 163 BUF1 $T=523900 739320 0 0 $X=523900 $Y=738940
X52 1422 2 1 1496 BUF1 $T=523900 860280 1 0 $X=523900 $Y=854860
X53 1282 2 1 1483 BUF1 $T=527000 809880 0 0 $X=527000 $Y=809500
X54 1483 2 1 1512 BUF1 $T=528860 830040 0 0 $X=528860 $Y=829660
X55 1512 2 1 1436 BUF1 $T=533820 840120 0 180 $X=531340 $Y=834700
X56 1468 2 1 1521 BUF1 $T=533820 759480 1 0 $X=533820 $Y=754060
X57 1468 2 1 1527 BUF1 $T=534440 769560 0 0 $X=534440 $Y=769180
X58 1512 2 1 1490 BUF1 $T=536920 840120 1 180 $X=534440 $Y=839740
X59 1483 2 1 1541 BUF1 $T=536300 809880 0 0 $X=536300 $Y=809500
X60 163 2 1 1561 BUF1 $T=548080 739320 0 180 $X=545600 $Y=733900
X61 1541 2 1 1562 BUF1 $T=546220 809880 0 0 $X=546220 $Y=809500
X62 1521 2 1 1537 BUF1 $T=550560 749400 1 0 $X=550560 $Y=743980
X63 1551 2 1 1579 BUF1 $T=550560 769560 1 0 $X=550560 $Y=764140
X64 1512 2 1 1606 BUF1 $T=553040 840120 0 0 $X=553040 $Y=839740
X65 1521 2 1 1635 BUF1 $T=553660 749400 1 0 $X=553660 $Y=743980
X66 1632 2 1 1602 BUF1 $T=558620 809880 0 0 $X=558620 $Y=809500
X67 1606 2 1 1622 BUF1 $T=559860 860280 1 0 $X=559860 $Y=854860
X68 1632 2 1 1595 BUF1 $T=564820 819960 1 180 $X=562340 $Y=819580
X69 1552 2 1 1660 BUF1 $T=562960 850200 1 0 $X=562960 $Y=844780
X70 1622 2 1 1661 BUF1 $T=563580 860280 0 0 $X=563580 $Y=859900
X71 1606 2 1 1668 BUF1 $T=566060 830040 0 0 $X=566060 $Y=829660
X72 175 2 1 1609 BUF1 $T=571640 890520 0 180 $X=569160 $Y=885100
X73 1635 2 1 1703 BUF1 $T=574120 749400 1 0 $X=574120 $Y=743980
X74 1659 2 1 1745 BUF1 $T=582180 749400 0 0 $X=582180 $Y=749020
X75 1750 2 1 1632 BUF1 $T=586520 819960 0 180 $X=584040 $Y=814540
X76 1660 2 1 1750 BUF1 $T=584040 850200 0 0 $X=584040 $Y=849820
X77 1728 2 1 184 BUF1 $T=587140 890520 1 180 $X=584660 $Y=890140
X78 1722 2 1 1680 BUF1 $T=586520 779640 0 0 $X=586520 $Y=779260
X79 1632 2 1 1762 BUF1 $T=587760 809880 0 0 $X=587760 $Y=809500
X80 1680 2 1 1781 BUF1 $T=589000 789720 0 0 $X=589000 $Y=789340
X81 1750 2 1 1772 BUF1 $T=589620 840120 0 0 $X=589620 $Y=839740
X82 1796 2 1 1728 BUF1 $T=592100 870360 1 0 $X=592100 $Y=864940
X83 1728 2 1 194 BUF1 $T=592100 890520 0 0 $X=592100 $Y=890140
X84 1722 2 1 1798 BUF1 $T=596440 759480 0 0 $X=596440 $Y=759100
X85 1790 2 1 1710 BUF1 $T=601400 799800 1 180 $X=598920 $Y=799420
X86 1776 2 1 1827 BUF1 $T=602020 830040 1 0 $X=602020 $Y=824620
X87 1798 2 1 1828 BUF1 $T=602640 769560 0 0 $X=602640 $Y=769180
X88 1772 2 1 1842 BUF1 $T=604500 850200 1 0 $X=604500 $Y=844780
X89 1837 2 1 1540 BUF1 $T=607600 759480 0 0 $X=607600 $Y=759100
X90 177 2 1 1682 BUF1 $T=611320 739320 1 0 $X=611320 $Y=733900
X91 1868 2 1 1776 BUF1 $T=611940 819960 1 0 $X=611940 $Y=814540
X92 1883 2 1 1790 BUF1 $T=618140 779640 1 180 $X=615660 $Y=779260
X93 1883 2 1 1868 BUF1 $T=620000 789720 0 180 $X=617520 $Y=784300
X94 1894 2 1 1322 BUF1 $T=618760 789720 0 0 $X=618760 $Y=789340
X95 1826 2 1 1909 BUF1 $T=621860 870360 0 0 $X=621860 $Y=869980
X96 1868 2 1 1917 BUF1 $T=623100 819960 1 0 $X=623100 $Y=814540
X97 1833 2 1 1932 BUF1 $T=624340 759480 0 0 $X=624340 $Y=759100
X98 1943 2 1 1894 BUF1 $T=628680 789720 0 0 $X=628680 $Y=789340
X99 1907 2 1 1938 BUF1 $T=630540 819960 1 0 $X=630540 $Y=814540
X100 1909 2 1 1920 BUF1 $T=634260 870360 1 180 $X=631780 $Y=869980
X101 1917 2 1 1921 BUF1 $T=634260 840120 1 0 $X=634260 $Y=834700
X102 1917 2 1 1955 BUF1 $T=637980 809880 0 180 $X=635500 $Y=804460
X103 231 2 1 1952 BUF1 $T=639220 890520 1 180 $X=636740 $Y=890140
X104 1982 2 1 1947 BUF1 $T=640460 840120 1 180 $X=637980 $Y=839740
X105 1980 2 1 1979 BUF1 $T=638600 759480 0 0 $X=638600 $Y=759100
X106 219 2 1 1999 BUF1 $T=639220 900600 1 0 $X=639220 $Y=895180
X107 1917 2 1 2000 BUF1 $T=639840 819960 0 0 $X=639840 $Y=819580
X108 1932 2 1 1883 BUF1 $T=641700 769560 0 0 $X=641700 $Y=769180
X109 1980 2 1 1906 BUF1 $T=642320 789720 1 0 $X=642320 $Y=784300
X110 1932 2 1 2049 BUF1 $T=649140 769560 0 0 $X=649140 $Y=769180
X111 231 2 1 2044 BUF1 $T=652240 890520 0 0 $X=652240 $Y=890140
X112 2006 2 1 2045 BUF1 $T=658440 749400 1 0 $X=658440 $Y=743980
X113 2096 2 1 254 BUF1 $T=665260 729240 0 0 $X=665260 $Y=728860
X114 2044 2 1 256 BUF1 $T=665260 900600 1 0 $X=665260 $Y=895180
X115 1982 2 1 2050 BUF1 $T=665880 840120 0 0 $X=665880 $Y=839740
X116 2044 2 1 2092 BUF1 $T=667740 890520 1 0 $X=667740 $Y=885100
X117 2012 2 1 2098 BUF1 $T=668980 789720 0 0 $X=668980 $Y=789340
X118 2050 2 1 2085 BUF1 $T=669600 830040 0 0 $X=669600 $Y=829660
X119 2043 2 1 2123 BUF1 $T=669600 860280 0 0 $X=669600 $Y=859900
X120 2043 2 1 2083 BUF1 $T=669600 880440 1 0 $X=669600 $Y=875020
X121 2153 2 1 2075 BUF1 $T=680760 799800 0 180 $X=678280 $Y=794380
X122 2085 2 1 2156 BUF1 $T=678900 819960 0 0 $X=678900 $Y=819580
X123 2107 2 1 2135 BUF1 $T=684480 759480 1 180 $X=682000 $Y=759100
X124 2135 2 1 2153 BUF1 $T=685720 789720 1 180 $X=683240 $Y=789340
X125 2083 2 1 2208 BUF1 $T=688200 890520 1 0 $X=688200 $Y=885100
X126 2085 2 1 2188 BUF1 $T=693780 830040 1 180 $X=691300 $Y=829660
X127 2208 2 1 274 BUF1 $T=696880 890520 1 180 $X=694400 $Y=890140
X128 2153 2 1 2209 BUF1 $T=696880 799800 1 0 $X=696880 $Y=794380
X129 283 2 1 2258 BUF1 $T=705560 729240 1 0 $X=705560 $Y=723820
X130 2247 2 1 2221 BUF1 $T=705560 870360 1 0 $X=705560 $Y=864940
X131 2200 2 1 292 BUF1 $T=707420 850200 0 0 $X=707420 $Y=849820
X132 2275 2 1 294 BUF1 $T=714240 900600 0 180 $X=711760 $Y=895180
X133 2208 2 1 2275 BUF1 $T=716720 890520 1 180 $X=714240 $Y=890140
X134 2235 2 1 2327 BUF1 $T=717960 739320 0 0 $X=717960 $Y=738940
X135 2280 2 1 2346 BUF1 $T=721680 840120 1 0 $X=721680 $Y=834700
X136 308 2 1 2247 BUF1 $T=725400 880440 1 180 $X=722920 $Y=880060
X137 308 2 1 2354 BUF1 $T=726020 880440 0 0 $X=726020 $Y=880060
X138 2370 2 1 2277 BUF1 $T=729740 779640 1 180 $X=727260 $Y=779260
X139 2280 2 1 2314 BUF1 $T=730360 819960 0 180 $X=727880 $Y=814540
X140 312 2 1 315 BUF1 $T=728500 739320 1 0 $X=728500 $Y=733900
X141 2275 2 1 316 BUF1 $T=728500 900600 1 0 $X=728500 $Y=895180
X142 2275 2 1 2300 BUF1 $T=729120 890520 0 0 $X=729120 $Y=890140
X143 298 2 1 2382 BUF1 $T=733460 759480 1 0 $X=733460 $Y=754060
X144 193 2 1 325 BUF1 $T=733460 799800 1 0 $X=733460 $Y=794380
X145 2346 2 1 2391 BUF1 $T=739660 840120 0 180 $X=737180 $Y=834700
X146 2346 2 1 2433 BUF1 $T=743380 819960 1 0 $X=743380 $Y=814540
X147 2433 2 1 2370 BUF1 $T=747720 789720 1 180 $X=745240 $Y=789340
X148 2346 2 1 2462 BUF1 $T=748960 840120 1 0 $X=748960 $Y=834700
X149 2487 2 1 2430 BUF1 $T=754540 819960 0 0 $X=754540 $Y=819580
X150 2553 2 1 2487 BUF1 $T=768180 819960 1 180 $X=765700 $Y=819580
X151 2462 2 1 2563 BUF1 $T=771900 840120 1 0 $X=771900 $Y=834700
X152 2589 2 1 357 BUF1 $T=774380 900600 0 180 $X=771900 $Y=895180
X153 220 2 1 2506 BUF1 $T=773760 870360 0 0 $X=773760 $Y=869980
X154 2506 2 1 2621 BUF1 $T=776240 860280 1 0 $X=776240 $Y=854860
X155 2474 2 1 2643 BUF1 $T=784300 799800 0 0 $X=784300 $Y=799420
X156 2643 2 1 2553 BUF1 $T=786780 819960 0 180 $X=784300 $Y=814540
X157 2648 2 1 2583 BUF1 $T=788020 880440 1 180 $X=785540 $Y=880060
X158 2621 2 1 2661 BUF1 $T=788020 819960 1 0 $X=788020 $Y=814540
X159 2589 2 1 369 BUF1 $T=788640 900600 1 0 $X=788640 $Y=895180
X160 2666 2 1 2589 BUF1 $T=791740 870360 1 180 $X=789260 $Y=869980
X161 2671 2 1 2601 BUF1 $T=792980 850200 1 180 $X=790500 $Y=849820
X162 2643 2 1 2680 BUF1 $T=796700 819960 0 180 $X=794220 $Y=814540
X163 2648 2 1 2671 BUF1 $T=795460 860280 1 0 $X=795460 $Y=854860
X164 2680 2 1 2666 BUF1 $T=796080 840120 0 0 $X=796080 $Y=839740
X165 2666 2 1 2716 BUF1 $T=799800 870360 0 0 $X=799800 $Y=869980
X166 2732 2 1 2728 BUF1 $T=804760 759480 0 0 $X=804760 $Y=759100
X167 2671 2 1 2755 BUF1 $T=812820 840120 1 0 $X=812820 $Y=834700
X168 2755 2 1 2749 BUF1 $T=819640 830040 0 180 $X=817160 $Y=824620
X169 393 2 1 392 BUF1 $T=817780 900600 1 0 $X=817780 $Y=895180
X170 2755 2 1 2800 BUF1 $T=820880 830040 1 0 $X=820880 $Y=824620
X171 2643 2 1 2832 BUF1 $T=823980 809880 1 0 $X=823980 $Y=804460
X172 2825 2 1 2732 BUF1 $T=830180 769560 0 180 $X=827700 $Y=764140
X173 2825 2 1 2873 BUF1 $T=839480 769560 0 180 $X=837000 $Y=764140
X174 2832 2 1 2811 BUF1 $T=840100 809880 1 0 $X=840100 $Y=804460
X175 2825 2 1 2902 BUF1 $T=841960 779640 1 0 $X=841960 $Y=774220
X176 2861 2 1 2825 BUF1 $T=845060 789720 1 180 $X=842580 $Y=789340
X177 2873 2 1 425 BUF1 $T=846920 749400 0 180 $X=844440 $Y=743980
X178 2851 2 1 2861 BUF1 $T=844440 809880 1 0 $X=844440 $Y=804460
X179 2811 2 1 3003 BUF1 $T=857460 799800 1 0 $X=857460 $Y=794380
X180 2932 2 1 3009 BUF1 $T=859320 870360 1 0 $X=859320 $Y=864940
X181 3001 2 1 3006 BUF1 $T=859940 789720 1 0 $X=859940 $Y=784300
X182 2851 2 1 3063 BUF1 $T=867380 819960 0 0 $X=867380 $Y=819580
X183 2920 2 1 3069 BUF1 $T=868000 759480 1 0 $X=868000 $Y=754060
X184 3146 2 1 3145 BUF1 $T=881020 759480 0 0 $X=881020 $Y=759100
X185 3114 2 1 3171 BUF1 $T=882880 840120 1 0 $X=882880 $Y=834700
X186 3063 2 1 3084 BUF1 $T=885980 819960 1 180 $X=883500 $Y=819580
X187 3009 2 1 3168 BUF1 $T=883500 870360 1 0 $X=883500 $Y=864940
X188 3063 2 1 3106 BUF1 $T=887220 809880 0 0 $X=887220 $Y=809500
X189 450 2 1 470 BUF1 $T=890940 890520 0 0 $X=890940 $Y=890140
X190 3083 2 1 3195 BUF1 $T=894660 749400 0 0 $X=894660 $Y=749020
X191 3063 2 1 3221 BUF1 $T=896520 809880 0 0 $X=896520 $Y=809500
X192 3245 2 1 481 BUF1 $T=899620 759480 1 0 $X=899620 $Y=754060
X193 3075 2 1 3280 BUF1 $T=903960 749400 0 0 $X=903960 $Y=749020
X194 3069 2 1 3307 BUF1 $T=906440 739320 1 0 $X=906440 $Y=733900
X195 3350 2 1 3353 BUF1 $T=916360 789720 0 0 $X=916360 $Y=789340
X196 3001 2 1 3343 BUF1 $T=923180 749400 0 0 $X=923180 $Y=749020
X197 3221 2 1 3425 BUF1 $T=930620 809880 0 0 $X=930620 $Y=809500
X198 3001 2 1 3488 BUF1 $T=940540 749400 0 0 $X=940540 $Y=749020
X199 3200 2 1 3521 BUF1 $T=946740 739320 0 0 $X=946740 $Y=738940
X200 3425 2 1 3420 BUF1 $T=956660 819960 1 0 $X=956660 $Y=814540
X201 3678 2 1 3661 BUF1 $T=1009360 719160 1 180 $X=1006880 $Y=718780
X202 3682 2 1 3664 BUF1 $T=1016180 769560 1 180 $X=1013700 $Y=769180
X203 3696 2 1 3682 BUF1 $T=1034160 769560 1 180 $X=1031680 $Y=769180
X204 3707 2 1 3710 BUF1 $T=1040360 749400 0 0 $X=1040360 $Y=749020
X205 3707 2 1 3722 BUF1 $T=1045320 749400 0 0 $X=1045320 $Y=749020
X206 3696 2 1 3712 BUF1 $T=1047180 769560 1 0 $X=1047180 $Y=764140
X207 567 2 1 3713 BUF1 $T=1058960 729240 0 180 $X=1056480 $Y=723820
X208 3712 2 1 3730 BUF1 $T=1056480 779640 1 0 $X=1056480 $Y=774220
X209 3697 2 1 3740 BUF1 $T=1062680 789720 0 0 $X=1062680 $Y=789340
X210 802 27 756 2 1 741 QDFFRBN $T=367660 890520 0 180 $X=355880 $Y=885100
X211 792 27 756 2 1 750 QDFFRBN $T=368280 880440 1 180 $X=356500 $Y=880060
X212 808 27 824 2 1 861 QDFFRBN $T=370140 860280 0 0 $X=370140 $Y=859900
X213 809 27 756 2 1 859 QDFFRBN $T=370140 890520 1 0 $X=370140 $Y=885100
X214 814 27 824 2 1 842 QDFFRBN $T=370760 870360 1 0 $X=370760 $Y=864940
X215 839 27 886 2 1 879 QDFFRBN $T=378200 860280 1 0 $X=378200 $Y=854860
X216 922 882 894 2 1 872 QDFFRBN $T=395560 830040 1 180 $X=383780 $Y=829660
X217 874 882 894 2 1 928 QDFFRBN $T=383780 840120 0 0 $X=383780 $Y=839740
X218 865 27 923 2 1 938 QDFFRBN $T=386260 880440 0 0 $X=386260 $Y=880060
X219 895 882 886 2 1 944 QDFFRBN $T=387500 850200 0 0 $X=387500 $Y=849820
X220 927 27 824 2 1 887 QDFFRBN $T=400520 870360 0 180 $X=388740 $Y=864940
X221 896 27 923 2 1 949 QDFFRBN $T=391840 890520 0 0 $X=391840 $Y=890140
X222 890 27 923 2 1 909 QDFFRBN $T=404240 890520 0 180 $X=392460 $Y=885100
X223 997 882 943 2 1 924 QDFFRBN $T=407340 819960 0 180 $X=395560 $Y=814540
X224 947 882 943 2 1 1000 QDFFRBN $T=399280 830040 0 0 $X=399280 $Y=829660
X225 956 882 886 2 1 1024 QDFFRBN $T=401760 860280 1 0 $X=401760 $Y=854860
X226 957 27 923 2 1 988 QDFFRBN $T=401760 880440 0 0 $X=401760 $Y=880060
X227 972 27 54 2 1 1026 QDFFRBN $T=404240 900600 1 0 $X=404240 $Y=895180
X228 995 27 1032 2 1 1043 QDFFRBN $T=408580 890520 1 0 $X=408580 $Y=885100
X229 1016 882 1029 2 1 1051 QDFFRBN $T=411680 830040 1 0 $X=411680 $Y=824620
X230 1057 882 1029 2 1 1004 QDFFRBN $T=424700 819960 0 180 $X=412920 $Y=814540
X231 1058 882 992 2 1 1019 QDFFRBN $T=425320 840120 1 180 $X=413540 $Y=839740
X232 1055 882 992 2 1 1023 QDFFRBN $T=425320 850200 0 180 $X=413540 $Y=844780
X233 1027 27 935 2 1 1068 QDFFRBN $T=415400 870360 1 0 $X=415400 $Y=864940
X234 71 27 1032 2 1 1100 QDFFRBN $T=422220 890520 0 0 $X=422220 $Y=890140
X235 1095 882 1070 2 1 1054 QDFFRBN $T=435240 799800 1 180 $X=423460 $Y=799420
X236 1096 882 1029 2 1 1036 QDFFRBN $T=435240 809880 1 180 $X=423460 $Y=809500
X237 1061 27 1032 2 1 1102 QDFFRBN $T=423460 880440 0 0 $X=423460 $Y=880060
X238 1104 882 1070 2 1 851 QDFFRBN $T=436480 799800 0 180 $X=424700 $Y=794380
X239 1064 882 1090 2 1 1105 QDFFRBN $T=424700 840120 1 0 $X=424700 $Y=834700
X240 1106 882 1070 2 1 834 QDFFRBN $T=437100 789720 1 180 $X=425320 $Y=789340
X241 1111 882 992 2 1 1066 QDFFRBN $T=437720 850200 0 180 $X=425940 $Y=844780
X242 1138 78 1097 2 1 1081 QDFFRBN $T=442680 860280 0 180 $X=430900 $Y=854860
X243 1084 78 1122 2 1 1139 QDFFRBN $T=430900 870360 1 0 $X=430900 $Y=864940
X244 1085 78 1122 2 1 1140 QDFFRBN $T=430900 880440 1 0 $X=430900 $Y=875020
X245 1136 882 1070 2 1 833 QDFFRBN $T=444540 789720 0 180 $X=432760 $Y=784300
X246 1107 78 87 2 1 1147 QDFFRBN $T=435240 890520 0 0 $X=435240 $Y=890140
X247 1118 882 1070 2 1 1155 QDFFRBN $T=437720 799800 1 0 $X=437720 $Y=794380
X248 1120 882 1090 2 1 1150 QDFFRBN $T=438960 840120 1 0 $X=438960 $Y=834700
X249 1166 78 1097 2 1 1121 QDFFRBN $T=450740 850200 1 180 $X=438960 $Y=849820
X250 1161 882 1131 2 1 829 QDFFRBN $T=451980 779640 1 180 $X=440200 $Y=779260
X251 1164 882 1131 2 1 845 QDFFRBN $T=453220 759480 1 180 $X=441440 $Y=759100
X252 1165 882 1131 2 1 827 QDFFRBN $T=453220 769560 0 180 $X=441440 $Y=764140
X253 1170 882 1131 2 1 831 QDFFRBN $T=453840 769560 1 180 $X=442060 $Y=769180
X254 1171 882 1131 2 1 841 QDFFRBN $T=453840 779640 0 180 $X=442060 $Y=774220
X255 1137 882 1133 2 1 1178 QDFFRBN $T=442680 819960 1 0 $X=442680 $Y=814540
X256 1141 882 1163 2 1 1180 QDFFRBN $T=443920 830040 0 0 $X=443920 $Y=829660
X257 1189 882 1133 2 1 1142 QDFFRBN $T=456320 809880 0 180 $X=444540 $Y=804460
X258 1144 78 1122 2 1 1159 QDFFRBN $T=445160 880440 1 0 $X=445160 $Y=875020
X259 1196 882 1133 2 1 1156 QDFFRBN $T=460040 809880 1 180 $X=448260 $Y=809500
X260 1199 6 953 2 1 1035 QDFFRBN $T=462520 739320 0 180 $X=450740 $Y=733900
X261 1200 6 953 2 1 973 QDFFRBN $T=462520 739320 1 180 $X=450740 $Y=738940
X262 1204 882 953 2 1 53 QDFFRBN $T=463140 749400 1 180 $X=451360 $Y=749020
X263 1205 882 953 2 1 91 QDFFRBN $T=463140 759480 0 180 $X=451360 $Y=754060
X264 107 78 100 2 1 1158 QDFFRBN $T=463140 890520 1 180 $X=451360 $Y=890140
X265 1192 882 1163 2 1 1169 QDFFRBN $T=465000 840120 1 180 $X=453220 $Y=839740
X266 1160 78 1122 2 1 1175 QDFFRBN $T=465000 860280 1 180 $X=453220 $Y=859900
X267 1193 78 1122 2 1 1173 QDFFRBN $T=465620 860280 0 180 $X=453840 $Y=854860
X268 1201 882 1154 2 1 1168 QDFFRBN $T=466240 789720 1 180 $X=454460 $Y=789340
X269 1233 78 1122 2 1 1181 QDFFRBN $T=466860 870360 1 180 $X=455080 $Y=869980
X270 1188 882 1154 2 1 1223 QDFFRBN $T=456320 769560 0 0 $X=456320 $Y=769180
X271 1225 882 1154 2 1 1179 QDFFRBN $T=468100 779640 0 180 $X=456320 $Y=774220
X272 1217 882 1163 2 1 1186 QDFFRBN $T=468100 840120 0 180 $X=456320 $Y=834700
X273 1219 882 1154 2 1 1182 QDFFRBN $T=468720 789720 0 180 $X=456940 $Y=784300
X274 1230 882 1133 2 1 1190 QDFFRBN $T=468720 809880 0 180 $X=456940 $Y=804460
X275 1198 882 1227 2 1 1231 QDFFRBN $T=460040 809880 0 0 $X=460040 $Y=809500
X276 1194 78 1234 2 1 1244 QDFFRBN $T=461280 890520 1 0 $X=461280 $Y=885100
X277 1218 78 100 2 1 105 QDFFRBN $T=473060 900600 0 180 $X=461280 $Y=895180
X278 1248 6 953 2 1 892 QDFFRBN $T=474300 749400 0 180 $X=462520 $Y=743980
X279 1167 78 1234 2 1 1207 QDFFRBN $T=462520 880440 0 0 $X=462520 $Y=880060
X280 1255 6 1220 2 1 982 QDFFRBN $T=476160 739320 1 180 $X=464380 $Y=738940
X281 1256 6 953 2 1 912 QDFFRBN $T=476160 749400 1 180 $X=464380 $Y=749020
X282 1212 882 1220 2 1 1261 QDFFRBN $T=464380 759480 0 0 $X=464380 $Y=759100
X283 1264 6 1220 2 1 1001 QDFFRBN $T=476780 739320 0 180 $X=465000 $Y=733900
X284 1208 882 1227 2 1 1202 QDFFRBN $T=465000 799800 0 0 $X=465000 $Y=799420
X285 1214 78 1250 2 1 1247 QDFFRBN $T=465620 850200 1 0 $X=465620 $Y=844780
X286 1221 78 1250 2 1 1268 QDFFRBN $T=466860 860280 1 0 $X=466860 $Y=854860
X287 1232 882 1250 2 1 1253 QDFFRBN $T=468720 840120 1 0 $X=468720 $Y=834700
X288 1237 882 1227 2 1 1289 QDFFRBN $T=469960 789720 0 0 $X=469960 $Y=789340
X289 1239 78 1234 2 1 1273 QDFFRBN $T=469960 870360 0 0 $X=469960 $Y=869980
X290 1243 6 122 2 1 1295 QDFFRBN $T=471200 729240 1 0 $X=471200 $Y=723820
X291 1290 882 1227 2 1 1242 QDFFRBN $T=482980 809880 0 180 $X=471200 $Y=804460
X292 1266 78 1234 2 1 1249 QDFFRBN $T=484840 890520 0 180 $X=473060 $Y=885100
X293 1252 882 1227 2 1 1311 QDFFRBN $T=473680 799800 1 0 $X=473680 $Y=794380
X294 1257 78 1234 2 1 1310 QDFFRBN $T=474300 900600 1 0 $X=474300 $Y=895180
X295 1263 882 1308 2 1 1323 QDFFRBN $T=476160 830040 1 0 $X=476160 $Y=824620
X296 1319 882 1286 2 1 1267 QDFFRBN $T=489180 759480 1 180 $X=477400 $Y=759100
X297 1269 882 1286 2 1 1324 QDFFRBN $T=477400 779640 1 0 $X=477400 $Y=774220
X298 1277 6 1220 2 1 1333 QDFFRBN $T=478640 739320 1 0 $X=478640 $Y=733900
X299 1291 78 1315 2 1 1341 QDFFRBN $T=481120 880440 0 0 $X=481120 $Y=880060
X300 1292 882 1286 2 1 1342 QDFFRBN $T=481740 769560 1 0 $X=481740 $Y=764140
X301 1284 882 1250 2 1 1340 QDFFRBN $T=481740 850200 0 0 $X=481740 $Y=849820
X302 1345 130 1315 2 1 1296 QDFFRBN $T=494140 870360 1 180 $X=482360 $Y=869980
X303 1347 1339 1308 2 1 1301 QDFFRBN $T=494760 809880 0 180 $X=482980 $Y=804460
X304 1298 882 1337 2 1 1283 QDFFRBN $T=482980 840120 1 0 $X=482980 $Y=834700
X305 1303 882 1337 2 1 1294 QDFFRBN $T=482980 850200 1 0 $X=482980 $Y=844780
X306 1304 882 1250 2 1 1348 QDFFRBN $T=482980 860280 1 0 $X=482980 $Y=854860
X307 1344 882 1308 2 1 1306 QDFFRBN $T=495380 819960 1 180 $X=483600 $Y=819580
X308 1317 6 122 2 1 1362 QDFFRBN $T=485460 729240 1 0 $X=485460 $Y=723820
X309 1320 78 1234 2 1 1361 QDFFRBN $T=486080 890520 0 0 $X=486080 $Y=890140
X310 1330 882 1360 2 1 1371 QDFFRBN $T=489180 799800 0 0 $X=489180 $Y=799420
X311 1328 78 139 2 1 1372 QDFFRBN $T=489180 900600 1 0 $X=489180 $Y=895180
X312 1334 882 1286 2 1 1375 QDFFRBN $T=490420 759480 0 0 $X=490420 $Y=759100
X313 1321 1339 1360 2 1 1389 QDFFRBN $T=492280 789720 0 0 $X=492280 $Y=789340
X314 1350 130 1315 2 1 1397 QDFFRBN $T=494140 880440 1 0 $X=494140 $Y=875020
X315 1352 882 1286 2 1 1380 QDFFRBN $T=494760 769560 1 0 $X=494760 $Y=764140
X316 1355 130 1315 2 1 1399 QDFFRBN $T=495380 870360 0 0 $X=495380 $Y=869980
X317 1363 1339 1368 2 1 1357 QDFFRBN $T=507780 850200 0 180 $X=496000 $Y=844780
X318 1394 130 1368 2 1 1354 QDFFRBN $T=508400 860280 0 180 $X=496620 $Y=854860
X319 1402 1339 1308 2 1 1377 QDFFRBN $T=513360 809880 1 180 $X=501580 $Y=809500
X320 1420 1339 1395 2 1 1378 QDFFRBN $T=513360 819960 1 180 $X=501580 $Y=819580
X321 142 133 149 2 1 153 QDFFRBN $T=502200 719160 0 0 $X=502200 $Y=718780
X322 1386 133 149 2 1 1428 QDFFRBN $T=502200 729240 1 0 $X=502200 $Y=723820
X323 1424 1339 1360 2 1 1383 QDFFRBN $T=513980 789720 0 180 $X=502200 $Y=784300
X324 1391 882 1286 2 1 1434 QDFFRBN $T=503440 759480 0 0 $X=503440 $Y=759100
X325 1404 1339 1360 2 1 1392 QDFFRBN $T=518320 799800 0 180 $X=506540 $Y=794380
X326 1405 1339 1422 2 1 1454 QDFFRBN $T=508400 850200 1 0 $X=508400 $Y=844780
X327 1410 1339 1447 2 1 1449 QDFFRBN $T=509640 840120 1 0 $X=509640 $Y=834700
X328 1411 130 1422 2 1 1466 QDFFRBN $T=509640 860280 1 0 $X=509640 $Y=854860
X329 1456 130 1422 2 1 1408 QDFFRBN $T=521420 870360 0 180 $X=509640 $Y=864940
X330 1425 1339 1447 2 1 1473 QDFFRBN $T=512120 830040 1 0 $X=512120 $Y=824620
X331 1471 1339 1414 2 1 1429 QDFFRBN $T=525140 789720 1 180 $X=513360 $Y=789340
X332 1433 1339 1414 2 1 1481 QDFFRBN $T=513980 789720 1 0 $X=513980 $Y=784300
X333 1407 1339 1468 2 1 1487 QDFFRBN $T=514600 779640 1 0 $X=514600 $Y=774220
X334 1441 1339 1458 2 1 1478 QDFFRBN $T=515220 809880 1 0 $X=515220 $Y=804460
X335 1482 1339 1395 2 1 1439 QDFFRBN $T=527000 819960 1 180 $X=515220 $Y=819580
X336 1440 133 149 2 1 166 QDFFRBN $T=519560 719160 0 0 $X=519560 $Y=718780
X337 1445 133 149 2 1 1469 QDFFRBN $T=519560 729240 1 0 $X=519560 $Y=723820
X338 1446 133 1468 2 1 1453 QDFFRBN $T=519560 759480 0 0 $X=519560 $Y=759100
X339 1442 130 1422 2 1 1500 QDFFRBN $T=520180 880440 1 0 $X=520180 $Y=875020
X340 1462 133 1468 2 1 1509 QDFFRBN $T=520800 759480 1 0 $X=520800 $Y=754060
X341 1465 1339 1489 2 1 1517 QDFFRBN $T=521420 840120 0 0 $X=521420 $Y=839740
X342 1472 130 1496 2 1 1513 QDFFRBN $T=523280 870360 1 0 $X=523280 $Y=864940
X343 1474 1339 1489 2 1 1525 QDFFRBN $T=523900 850200 0 0 $X=523900 $Y=849820
X344 1484 130 168 2 1 1518 QDFFRBN $T=525140 900600 1 0 $X=525140 $Y=895180
X345 1475 130 1496 2 1 1531 QDFFRBN $T=525760 870360 0 0 $X=525760 $Y=869980
X346 1461 133 1521 2 1 1532 QDFFRBN $T=526380 749400 1 0 $X=526380 $Y=743980
X347 1467 130 168 2 1 1533 QDFFRBN $T=526380 890520 1 0 $X=526380 $Y=885100
X348 1495 1339 1468 2 1 1542 QDFFRBN $T=528240 779640 1 0 $X=528240 $Y=774220
X349 1519 1339 1458 2 1 1492 QDFFRBN $T=540020 799800 1 180 $X=528240 $Y=799420
X350 1511 1339 1458 2 1 1493 QDFFRBN $T=540020 809880 0 180 $X=528240 $Y=804460
X351 1501 133 1521 2 1 1559 QDFFRBN $T=529480 749400 0 0 $X=529480 $Y=749020
X352 1505 1339 1496 2 1 1555 QDFFRBN $T=530100 860280 1 0 $X=530100 $Y=854860
X353 1486 133 1537 2 1 1548 QDFFRBN $T=530720 729240 0 0 $X=530720 $Y=728860
X354 1545 130 168 2 1 1506 QDFFRBN $T=542500 880440 1 180 $X=530720 $Y=880060
X355 171 133 149 2 1 1507 QDFFRBN $T=543120 719160 1 180 $X=531340 $Y=718780
X356 1508 133 1537 2 1 1557 QDFFRBN $T=531340 739320 0 0 $X=531340 $Y=738940
X357 1516 1339 1447 2 1 1568 QDFFRBN $T=533200 830040 0 0 $X=533200 $Y=829660
X358 1563 1339 1447 2 1 1522 QDFFRBN $T=546220 819960 0 180 $X=534440 $Y=814540
X359 1523 1339 1447 2 1 1515 QDFFRBN $T=546220 830040 0 180 $X=534440 $Y=824620
X360 1524 1339 1496 2 1 1573 QDFFRBN $T=534440 850200 1 0 $X=534440 $Y=844780
X361 1575 1339 1527 2 1 1534 QDFFRBN $T=549940 769560 1 180 $X=538160 $Y=769180
X362 1558 133 1521 2 1 1603 QDFFRBN $T=542500 749400 0 0 $X=542500 $Y=749020
X363 1554 1339 1595 2 1 1605 QDFFRBN $T=543120 809880 1 0 $X=543120 $Y=804460
X364 1560 130 175 2 1 1588 QDFFRBN $T=543740 890520 0 0 $X=543740 $Y=890140
X365 1569 133 1537 2 1 1611 QDFFRBN $T=544360 739320 0 0 $X=544360 $Y=738940
X366 1570 130 1552 2 1 1601 QDFFRBN $T=544980 860280 1 0 $X=544980 $Y=854860
X367 1571 1339 1602 2 1 1616 QDFFRBN $T=545600 799800 0 0 $X=545600 $Y=799420
X368 1576 1339 1595 2 1 1614 QDFFRBN $T=545600 819960 0 0 $X=545600 $Y=819580
X369 1564 130 1496 2 1 1578 QDFFRBN $T=558000 850200 0 180 $X=546220 $Y=844780
X370 1580 130 1552 2 1 1630 QDFFRBN $T=546220 870360 1 0 $X=546220 $Y=864940
X371 1620 133 1521 2 1 1581 QDFFRBN $T=558620 759480 0 180 $X=546840 $Y=754060
X372 1618 1339 1527 2 1 1591 QDFFRBN $T=562340 769560 1 180 $X=550560 $Y=769180
X373 1597 130 1609 2 1 1663 QDFFRBN $T=555520 890520 1 0 $X=555520 $Y=885100
X374 1613 1339 1595 2 1 1672 QDFFRBN $T=556140 819960 1 0 $X=556140 $Y=814540
X375 1648 1339 1527 2 1 1612 QDFFRBN $T=568540 779640 0 180 $X=556760 $Y=774220
X376 1621 1339 1595 2 1 1655 QDFFRBN $T=556760 840120 1 0 $X=556760 $Y=834700
X377 1600 130 1552 2 1 1645 QDFFRBN $T=556760 850200 0 0 $X=556760 $Y=849820
X378 1626 1339 1595 2 1 1676 QDFFRBN $T=557380 830040 1 0 $X=557380 $Y=824620
X379 1629 1339 1602 2 1 1675 QDFFRBN $T=558000 809880 1 0 $X=558000 $Y=804460
X380 1633 130 175 2 1 1681 QDFFRBN $T=558620 890520 0 0 $X=558620 $Y=890140
X381 1636 130 1552 2 1 1677 QDFFRBN $T=559240 870360 1 0 $X=559240 $Y=864940
X382 1671 133 1635 2 1 1631 QDFFRBN $T=572260 759480 0 180 $X=560480 $Y=754060
X383 1642 133 1635 2 1 1687 QDFFRBN $T=561100 749400 1 0 $X=561100 $Y=743980
X384 1643 1339 1680 2 1 1634 QDFFRBN $T=561720 789720 0 0 $X=561720 $Y=789340
X385 1650 1339 1602 2 1 1693 QDFFRBN $T=564200 799800 0 0 $X=564200 $Y=799420
X386 1652 130 1660 2 1 1724 QDFFRBN $T=569780 850200 0 0 $X=569780 $Y=849820
X387 1674 130 185 2 1 1706 QDFFRBN $T=570400 880440 0 0 $X=570400 $Y=880060
X388 1707 130 175 2 1 1685 QDFFRBN $T=582180 890520 1 180 $X=570400 $Y=890140
X389 1686 133 1703 2 1 1737 QDFFRBN $T=571020 729240 1 0 $X=571020 $Y=723820
X390 1688 1339 1722 2 1 1683 QDFFRBN $T=571020 769560 1 0 $X=571020 $Y=764140
X391 1689 1339 1722 2 1 1739 QDFFRBN $T=571020 769560 0 0 $X=571020 $Y=769180
X392 1730 1733 1703 2 1 1695 QDFFRBN $T=584040 739320 1 180 $X=572260 $Y=738940
X393 1697 133 1635 2 1 1741 QDFFRBN $T=572260 759480 1 0 $X=572260 $Y=754060
X394 1694 130 1660 2 1 1742 QDFFRBN $T=572260 870360 1 0 $X=572260 $Y=864940
X395 1699 1339 1680 2 1 1753 QDFFRBN $T=574740 789720 0 0 $X=574740 $Y=789340
X396 1715 130 1751 2 1 1757 QDFFRBN $T=577220 880440 1 0 $X=577220 $Y=875020
X397 1718 130 1750 2 1 1768 QDFFRBN $T=577840 860280 0 0 $X=577840 $Y=859900
X398 1727 1339 1762 2 1 1770 QDFFRBN $T=579700 799800 0 0 $X=579700 $Y=799420
X399 1759 1733 1703 2 1 1725 QDFFRBN $T=592100 749400 0 180 $X=580320 $Y=743980
X400 1705 1339 1762 2 1 1777 QDFFRBN $T=580320 809880 1 0 $X=580320 $Y=804460
X401 1734 1339 1722 2 1 1764 QDFFRBN $T=580940 759480 0 0 $X=580940 $Y=759100
X402 1723 1339 1750 2 1 1786 QDFFRBN $T=583420 840120 1 0 $X=583420 $Y=834700
X403 188 130 185 2 1 195 QDFFRBN $T=583420 900600 1 0 $X=583420 $Y=895180
X404 1740 192 196 2 1 200 QDFFRBN $T=587140 719160 0 0 $X=587140 $Y=718780
X405 1799 1733 1703 2 1 1758 QDFFRBN $T=599540 729240 1 180 $X=587760 $Y=728860
X406 1793 198 1772 2 1 1763 QDFFRBN $T=599540 850200 1 180 $X=587760 $Y=849820
X407 1752 1339 1722 2 1 1805 QDFFRBN $T=589000 779640 0 0 $X=589000 $Y=779260
X408 1749 1733 1798 2 1 1816 QDFFRBN $T=589620 769560 0 0 $X=589620 $Y=769180
X409 1778 1733 1703 2 1 1821 QDFFRBN $T=591480 739320 1 0 $X=591480 $Y=733900
X410 1780 130 1751 2 1 1815 QDFFRBN $T=592100 880440 1 0 $X=592100 $Y=875020
X411 1784 1339 1762 2 1 1835 QDFFRBN $T=593960 809880 1 0 $X=593960 $Y=804460
X412 1792 1339 1772 2 1 1850 QDFFRBN $T=595820 840120 0 0 $X=595820 $Y=839740
X413 1851 1733 1798 2 1 1807 QDFFRBN $T=611320 769560 0 180 $X=599540 $Y=764140
X414 1787 198 1842 2 1 1866 QDFFRBN $T=600780 860280 0 0 $X=600780 $Y=859900
X415 1817 198 1842 2 1 1861 QDFFRBN $T=601400 870360 0 0 $X=601400 $Y=869980
X416 1814 1733 1828 2 1 1849 QDFFRBN $T=602020 779640 0 0 $X=602020 $Y=779260
X417 1859 1733 1762 2 1 1820 QDFFRBN $T=613800 799800 1 180 $X=602020 $Y=799420
X418 1825 1733 1863 2 1 1875 QDFFRBN $T=603260 749400 1 0 $X=603260 $Y=743980
X419 1802 1733 1781 2 1 1829 QDFFRBN $T=616900 789720 0 180 $X=605120 $Y=784300
X420 1818 198 1751 2 1 1890 QDFFRBN $T=605120 880440 1 0 $X=605120 $Y=875020
X421 1839 192 207 2 1 1877 QDFFRBN $T=605740 729240 1 0 $X=605740 $Y=723820
X422 1881 1733 1781 2 1 1838 QDFFRBN $T=617520 789720 1 180 $X=605740 $Y=789340
X423 1834 198 1751 2 1 1843 QDFFRBN $T=605740 880440 0 0 $X=605740 $Y=880060
X424 1884 1733 1762 2 1 1848 QDFFRBN $T=619380 809880 1 180 $X=607600 $Y=809500
X425 1852 1733 1828 2 1 1898 QDFFRBN $T=608840 779640 1 0 $X=608840 $Y=774220
X426 1853 198 1751 2 1 1905 QDFFRBN $T=608840 890520 0 0 $X=608840 $Y=890140
X427 1856 1733 1772 2 1 1903 QDFFRBN $T=609460 830040 0 0 $X=609460 $Y=829660
X428 1857 198 1772 2 1 1902 QDFFRBN $T=609460 840120 0 0 $X=609460 $Y=839740
X429 1864 198 1842 2 1 1896 QDFFRBN $T=611320 870360 1 0 $X=611320 $Y=864940
X430 1867 192 207 2 1 1916 QDFFRBN $T=611940 719160 0 0 $X=611940 $Y=718780
X431 1871 1733 1828 2 1 1908 QDFFRBN $T=612560 769560 0 0 $X=612560 $Y=769180
X432 1858 198 1842 2 1 1919 QDFFRBN $T=613180 860280 1 0 $X=613180 $Y=854860
X433 1874 1733 1906 2 1 1888 QDFFRBN $T=613800 799800 1 0 $X=613800 $Y=794380
X434 1872 1733 1907 2 1 1924 QDFFRBN $T=613800 830040 1 0 $X=613800 $Y=824620
X435 1910 1733 1863 2 1 1882 QDFFRBN $T=628060 749400 0 180 $X=616280 $Y=743980
X436 1889 1733 1863 2 1 1935 QDFFRBN $T=617520 739320 0 0 $X=617520 $Y=738940
X437 1944 1733 1863 2 1 1891 QDFFRBN $T=630540 759480 0 180 $X=618760 $Y=754060
X438 1904 1733 1938 2 1 1936 QDFFRBN $T=620620 809880 0 0 $X=620620 $Y=809500
X439 1911 198 1947 2 1 1959 QDFFRBN $T=622480 840120 0 0 $X=622480 $Y=839740
X440 1918 198 1952 2 1 1960 QDFFRBN $T=623720 890520 0 0 $X=623720 $Y=890140
X441 1922 198 1952 2 1 1965 QDFFRBN $T=624340 870360 1 0 $X=624340 $Y=864940
X442 1925 192 223 2 1 228 QDFFRBN $T=624960 719160 0 0 $X=624960 $Y=718780
X443 1926 1733 1906 2 1 1963 QDFFRBN $T=624960 779640 1 0 $X=624960 $Y=774220
X444 1901 198 1952 2 1 1968 QDFFRBN $T=624960 880440 1 0 $X=624960 $Y=875020
X445 1966 1733 1907 2 1 1927 QDFFRBN $T=637360 830040 0 180 $X=625580 $Y=824620
X446 1931 198 1907 2 1 1973 QDFFRBN $T=625580 830040 0 0 $X=625580 $Y=829660
X447 1946 1733 1906 2 1 1934 QDFFRBN $T=638600 799800 0 180 $X=626820 $Y=794380
X448 1939 1733 1906 2 1 1969 QDFFRBN $T=628680 789720 1 0 $X=628680 $Y=784300
X449 1940 198 1947 2 1 1988 QDFFRBN $T=628680 850200 1 0 $X=628680 $Y=844780
X450 1948 1733 1863 2 1 1977 QDFFRBN $T=630540 739320 0 0 $X=630540 $Y=738940
X451 1953 1733 1980 2 1 2002 QDFFRBN $T=631780 769560 1 0 $X=631780 $Y=764140
X452 1957 198 1951 2 1 2011 QDFFRBN $T=633020 860280 1 0 $X=633020 $Y=854860
X453 1958 1733 1938 2 1 2003 QDFFRBN $T=633640 809880 0 0 $X=633640 $Y=809500
X454 1971 1733 1956 2 1 2022 QDFFRBN $T=636740 729240 0 0 $X=636740 $Y=728860
X455 1972 1733 1906 2 1 2018 QDFFRBN $T=636740 789720 0 0 $X=636740 $Y=789340
X456 1978 1733 1906 2 1 2026 QDFFRBN $T=637980 779640 1 0 $X=637980 $Y=774220
X457 1983 198 1952 2 1 2034 QDFFRBN $T=638600 880440 1 0 $X=638600 $Y=875020
X458 2024 192 1956 2 1 1987 QDFFRBN $T=651620 739320 0 180 $X=639840 $Y=733900
X459 1993 1733 1907 2 1 2039 QDFFRBN $T=641080 819960 1 0 $X=641080 $Y=814540
X460 2020 198 1951 2 1 1997 QDFFRBN $T=654720 860280 1 180 $X=642940 $Y=859900
X461 1981 198 1982 2 1 2053 QDFFRBN $T=644800 840120 1 0 $X=644800 $Y=834700
X462 2013 1733 1980 2 1 2054 QDFFRBN $T=645420 789720 1 0 $X=645420 $Y=784300
X463 2015 198 1982 2 1 2058 QDFFRBN $T=646040 850200 0 0 $X=646040 $Y=849820
X464 2007 198 2044 2 1 2037 QDFFRBN $T=646040 890520 1 0 $X=646040 $Y=885100
X465 2060 1733 2012 2 1 2019 QDFFRBN $T=659680 809880 0 180 $X=647900 $Y=804460
X466 2025 192 1956 2 1 2072 QDFFRBN $T=649760 739320 0 0 $X=649760 $Y=738940
X467 2031 192 1956 2 1 2073 QDFFRBN $T=650380 729240 0 0 $X=650380 $Y=728860
X468 2069 1733 1980 2 1 2028 QDFFRBN $T=662160 779640 0 180 $X=650380 $Y=774220
X469 2071 198 2044 2 1 2030 QDFFRBN $T=662160 880440 1 180 $X=650380 $Y=880060
X470 2033 1733 2063 2 1 2027 QDFFRBN $T=651000 759480 0 0 $X=651000 $Y=759100
X471 2038 1733 2063 2 1 2081 QDFFRBN $T=651620 749400 0 0 $X=651620 $Y=749020
X472 2055 198 2078 2 1 2108 QDFFRBN $T=655960 860280 0 0 $X=655960 $Y=859900
X473 2114 1733 2012 2 1 2065 QDFFRBN $T=671460 799800 0 180 $X=659680 $Y=794380
X474 2067 1733 2012 2 1 2101 QDFFRBN $T=659680 809880 1 0 $X=659680 $Y=804460
X475 2070 198 2050 2 1 2128 QDFFRBN $T=660300 840120 1 0 $X=660300 $Y=834700
X476 2074 1733 2063 2 1 2088 QDFFRBN $T=660920 769560 1 0 $X=660920 $Y=764140
X477 2082 192 2096 2 1 2136 QDFFRBN $T=662780 739320 0 0 $X=662780 $Y=738940
X478 2117 2127 254 2 1 2084 QDFFRBN $T=675180 729240 0 180 $X=663400 $Y=723820
X479 2120 1733 2063 2 1 2090 QDFFRBN $T=676420 759480 0 180 $X=664640 $Y=754060
X480 2133 198 2078 2 1 2103 QDFFRBN $T=679520 850200 1 180 $X=667740 $Y=849820
X481 266 198 256 2 1 2104 QDFFRBN $T=679520 900600 0 180 $X=667740 $Y=895180
X482 2160 198 2092 2 1 2109 QDFFRBN $T=680760 880440 1 180 $X=668980 $Y=880060
X483 2113 1733 2147 2 1 2162 QDFFRBN $T=669600 769560 0 0 $X=669600 $Y=769180
X484 2100 1733 2085 2 1 2167 QDFFRBN $T=670840 830040 1 0 $X=670840 $Y=824620
X485 2174 198 2092 2 1 2116 QDFFRBN $T=682620 890520 1 180 $X=670840 $Y=890140
X486 2121 1733 2098 2 1 2148 QDFFRBN $T=671460 789720 0 0 $X=671460 $Y=789340
X487 2151 1733 2063 2 1 2130 QDFFRBN $T=684480 749400 1 180 $X=672700 $Y=749020
X488 2134 1733 2156 2 1 2182 QDFFRBN $T=673320 809880 0 0 $X=673320 $Y=809500
X489 2142 2127 2096 2 1 2195 QDFFRBN $T=675800 729240 0 0 $X=675800 $Y=728860
X490 2194 2127 2096 2 1 2140 QDFFRBN $T=687580 739320 1 180 $X=675800 $Y=738940
X491 2138 198 2078 2 1 2189 QDFFRBN $T=675800 870360 1 0 $X=675800 $Y=864940
X492 2145 198 2078 2 1 2192 QDFFRBN $T=676420 870360 0 0 $X=676420 $Y=869980
X493 2137 192 275 2 1 2142 QDFFRBN $T=678900 719160 0 0 $X=678900 $Y=718780
X494 2154 198 2188 2 1 2146 QDFFRBN $T=678900 840120 1 0 $X=678900 $Y=834700
X495 2131 198 2085 2 1 2216 QDFFRBN $T=679520 830040 0 0 $X=679520 $Y=829660
X496 2159 198 2188 2 1 2206 QDFFRBN $T=680140 850200 1 0 $X=680140 $Y=844780
X497 2152 2127 2096 2 1 2211 QDFFRBN $T=681380 739320 1 0 $X=681380 $Y=733900
X498 2165 2127 2156 2 1 2191 QDFFRBN $T=682620 819960 0 0 $X=682620 $Y=819580
X499 2173 270 2201 2 1 2215 QDFFRBN $T=682620 890520 0 0 $X=682620 $Y=890140
X500 2179 1733 2098 2 1 2213 QDFFRBN $T=684480 789720 1 0 $X=684480 $Y=784300
X501 2176 2127 2147 2 1 2223 QDFFRBN $T=685100 769560 0 0 $X=685100 $Y=769180
X502 2184 1733 2219 2 1 2212 QDFFRBN $T=686340 749400 0 0 $X=686340 $Y=749020
X503 2187 270 2201 2 1 2228 QDFFRBN $T=686340 880440 0 0 $X=686340 $Y=880060
X504 2190 2127 2156 2 1 2229 QDFFRBN $T=686960 809880 1 0 $X=686960 $Y=804460
X505 2166 270 2221 2 1 2233 QDFFRBN $T=687580 860280 0 0 $X=687580 $Y=859900
X506 276 270 2201 2 1 284 QDFFRBN $T=688200 900600 1 0 $X=688200 $Y=895180
X507 2197 2127 2156 2 1 2239 QDFFRBN $T=688820 819960 1 0 $X=688820 $Y=814540
X508 2198 270 2221 2 1 2232 QDFFRBN $T=688820 870360 1 0 $X=688820 $Y=864940
X509 2205 2127 2156 2 1 2253 QDFFRBN $T=690680 830040 1 0 $X=690680 $Y=824620
X510 2207 270 2221 2 1 2246 QDFFRBN $T=690680 860280 1 0 $X=690680 $Y=854860
X511 2211 2127 2219 2 1 289 QDFFRBN $T=692540 739320 0 0 $X=692540 $Y=738940
X512 2204 2127 2219 2 1 288 QDFFRBN $T=692540 749400 1 0 $X=692540 $Y=743980
X513 2212 2127 2219 2 1 2282 QDFFRBN $T=692540 759480 1 0 $X=692540 $Y=754060
X514 2218 2127 2243 2 1 2261 QDFFRBN $T=693780 779640 0 0 $X=693780 $Y=779260
X515 2272 270 2247 2 1 2225 QDFFRBN $T=710520 880440 0 180 $X=698740 $Y=875020
X516 2237 270 2221 2 1 2287 QDFFRBN $T=699360 870360 0 0 $X=699360 $Y=869980
X517 293 270 2201 2 1 285 QDFFRBN $T=711760 900600 0 180 $X=699980 $Y=895180
X518 286 2127 2243 2 1 296 QDFFRBN $T=700600 749400 0 0 $X=700600 $Y=749020
X519 2286 270 2201 2 1 2241 QDFFRBN $T=712380 890520 1 180 $X=700600 $Y=890140
X520 2245 270 2221 2 1 2296 QDFFRBN $T=701220 860280 0 0 $X=701220 $Y=859900
X521 2248 2127 2243 2 1 299 QDFFRBN $T=701840 759480 0 0 $X=701840 $Y=759100
X522 2249 2127 2277 2 1 2263 QDFFRBN $T=701840 779640 1 0 $X=701840 $Y=774220
X523 2252 2127 2243 2 1 2302 QDFFRBN $T=702460 789720 1 0 $X=702460 $Y=784300
X524 2255 2127 2280 2 1 2304 QDFFRBN $T=702460 840120 0 0 $X=702460 $Y=839740
X525 2260 2127 2280 2 1 2309 QDFFRBN $T=704320 830040 1 0 $X=704320 $Y=824620
X526 2254 2127 2280 2 1 2310 QDFFRBN $T=704320 830040 0 0 $X=704320 $Y=829660
X527 2250 2127 2243 2 1 2276 QDFFRBN $T=705560 769560 0 0 $X=705560 $Y=769180
X528 2238 2127 2243 2 1 2313 QDFFRBN $T=706180 769560 1 0 $X=706180 $Y=764140
X529 2270 2127 2314 2 1 2325 QDFFRBN $T=708040 819960 1 0 $X=708040 $Y=814540
X530 2293 2127 2277 2 1 311 QDFFRBN $T=712380 779640 0 0 $X=712380 $Y=779260
X531 2315 2127 2277 2 1 313 QDFFRBN $T=716100 779640 1 0 $X=716100 $Y=774220
X532 2279 2127 2346 2 1 2326 QDFFRBN $T=716100 840120 0 0 $X=716100 $Y=839740
X533 2317 270 308 2 1 2358 QDFFRBN $T=716720 890520 1 0 $X=716720 $Y=885100
X534 2284 2127 2314 2 1 2361 QDFFRBN $T=717340 809880 1 0 $X=717340 $Y=804460
X535 2291 270 2247 2 1 2372 QDFFRBN $T=718580 870360 1 0 $X=718580 $Y=864940
X536 2332 2127 2277 2 1 320 QDFFRBN $T=720440 769560 0 0 $X=720440 $Y=769180
X537 2340 2127 2370 2 1 321 QDFFRBN $T=722300 789720 1 0 $X=722300 $Y=784300
X538 2341 2127 2346 2 1 2352 QDFFRBN $T=722300 819960 0 0 $X=722300 $Y=819580
X539 2342 2127 2280 2 1 2390 QDFFRBN $T=724160 840120 1 0 $X=724160 $Y=834700
X540 2357 2127 2370 2 1 317 QDFFRBN $T=742760 789720 1 180 $X=730980 $Y=789340
X541 2398 270 308 2 1 2371 QDFFRBN $T=742760 880440 1 180 $X=730980 $Y=880060
X542 2381 2127 2370 2 1 334 QDFFRBN $T=732840 779640 0 0 $X=732840 $Y=779260
X543 2425 270 2354 2 1 2384 QDFFRBN $T=745860 880440 0 180 $X=734080 $Y=875020
X544 2394 2127 2346 2 1 2452 QDFFRBN $T=735320 819960 0 0 $X=735320 $Y=819580
X545 2453 270 308 2 1 2392 QDFFRBN $T=747100 890520 0 180 $X=735320 $Y=885100
X546 2388 2127 2370 2 1 343 QDFFRBN $T=735940 789720 1 0 $X=735940 $Y=784300
X547 2404 2127 2433 2 1 2457 QDFFRBN $T=737800 799800 1 0 $X=737800 $Y=794380
X548 2411 2127 2391 2 1 2466 QDFFRBN $T=740280 850200 1 0 $X=740280 $Y=844780
X549 2418 2127 2462 2 1 2468 QDFFRBN $T=741520 830040 0 0 $X=741520 $Y=829660
X550 2431 270 2391 2 1 2488 QDFFRBN $T=744000 860280 1 0 $X=744000 $Y=854860
X551 2440 270 338 2 1 2501 QDFFRBN $T=745860 880440 1 0 $X=745860 $Y=875020
X552 2448 270 338 2 1 347 QDFFRBN $T=747100 900600 1 0 $X=747100 $Y=895180
X553 2455 2127 2433 2 1 2517 QDFFRBN $T=748340 819960 1 0 $X=748340 $Y=814540
X554 2460 270 338 2 1 2518 QDFFRBN $T=748960 890520 1 0 $X=748960 $Y=885100
X555 2484 2127 2479 2 1 2542 QDFFRBN $T=753920 799800 0 0 $X=753920 $Y=799420
X556 2486 2127 2479 2 1 2543 QDFFRBN $T=754540 789720 0 0 $X=754540 $Y=789340
X557 2480 2127 2462 2 1 2510 QDFFRBN $T=754540 830040 0 0 $X=754540 $Y=829660
X558 2475 2127 2462 2 1 2565 QDFFRBN $T=757640 840120 1 0 $X=757640 $Y=834700
X559 2515 2127 2563 2 1 2577 QDFFRBN $T=759500 830040 1 0 $X=759500 $Y=824620
X560 2532 2127 2563 2 1 2582 QDFFRBN $T=762600 819960 1 0 $X=762600 $Y=814540
X561 2552 2127 2479 2 1 2606 QDFFRBN $T=766320 799800 1 0 $X=766320 $Y=794380
X562 2556 270 2583 2 1 2608 QDFFRBN $T=766320 890520 1 0 $X=766320 $Y=885100
X563 2566 270 2601 2 1 2617 QDFFRBN $T=768180 860280 0 0 $X=768180 $Y=859900
X564 2574 2127 2462 2 1 2623 QDFFRBN $T=770040 840120 0 0 $X=770040 $Y=839740
X565 2618 360 2479 2 1 2576 QDFFRBN $T=782440 789720 1 180 $X=770660 $Y=789340
X566 2555 2127 2601 2 1 2637 QDFFRBN $T=772520 850200 0 0 $X=772520 $Y=849820
X567 2602 270 364 2 1 366 QDFFRBN $T=775620 900600 1 0 $X=775620 $Y=895180
X568 2616 270 2583 2 1 2668 QDFFRBN $T=779340 890520 1 0 $X=779340 $Y=885100
X569 2615 2127 2563 2 1 2657 QDFFRBN $T=779960 830040 0 0 $X=779960 $Y=829660
X570 2622 2127 2563 2 1 2654 QDFFRBN $T=780580 840120 1 0 $X=780580 $Y=834700
X571 2636 360 2628 2 1 2683 QDFFRBN $T=783680 779640 0 0 $X=783680 $Y=779260
X572 365 360 2628 2 1 2685 QDFFRBN $T=784300 789720 1 0 $X=784300 $Y=784300
X573 2498 360 2628 2 1 2696 QDFFRBN $T=784300 789720 0 0 $X=784300 $Y=789340
X574 2642 360 2628 2 1 2684 QDFFRBN $T=784920 799800 1 0 $X=784920 $Y=794380
X575 2652 270 2648 2 1 2698 QDFFRBN $T=786780 860280 0 0 $X=786780 $Y=859900
X576 2653 270 2648 2 1 2699 QDFFRBN $T=786780 880440 1 0 $X=786780 $Y=875020
X577 2655 270 2601 2 1 2688 QDFFRBN $T=788020 850200 1 0 $X=788020 $Y=844780
X578 2677 270 2648 2 1 2726 QDFFRBN $T=792360 880440 0 0 $X=792360 $Y=880060
X579 2682 2687 2671 2 1 2737 QDFFRBN $T=794220 840120 1 0 $X=794220 $Y=834700
X580 2578 360 2628 2 1 2745 QDFFRBN $T=794840 779640 1 0 $X=794840 $Y=774220
X581 2670 360 2732 2 1 2743 QDFFRBN $T=797320 769560 0 0 $X=797320 $Y=769180
X582 2715 270 2671 2 1 2703 QDFFRBN $T=810340 860280 0 180 $X=798560 $Y=854860
X583 2697 2687 2747 2 1 2753 QDFFRBN $T=802280 809880 0 0 $X=802280 $Y=809500
X584 2714 270 2671 2 1 2754 QDFFRBN $T=802280 850200 1 0 $X=802280 $Y=844780
X585 2702 270 2671 2 1 2757 QDFFRBN $T=804140 850200 0 0 $X=804140 $Y=849820
X586 2707 2687 2755 2 1 2734 QDFFRBN $T=806000 830040 0 0 $X=806000 $Y=829660
X587 2723 360 2728 2 1 2770 QDFFRBN $T=807860 759480 1 0 $X=807860 $Y=754060
X588 2588 360 2728 2 1 2771 QDFFRBN $T=807860 759480 0 0 $X=807860 $Y=759100
X589 2597 360 2732 2 1 2783 QDFFRBN $T=807860 769560 1 0 $X=807860 $Y=764140
X590 2739 270 392 2 1 2752 QDFFRBN $T=807860 890520 1 0 $X=807860 $Y=885100
X591 2541 270 393 2 1 398 QDFFRBN $T=807860 890520 0 0 $X=807860 $Y=890140
X592 2691 2687 2747 2 1 2798 QDFFRBN $T=809100 799800 1 0 $X=809100 $Y=794380
X593 2740 270 392 2 1 2778 QDFFRBN $T=809720 860280 0 0 $X=809720 $Y=859900
X594 2736 270 392 2 1 2785 QDFFRBN $T=809720 880440 1 0 $X=809720 $Y=875020
X595 2733 270 392 2 1 2759 QDFFRBN $T=810340 870360 0 0 $X=810340 $Y=869980
X596 2791 360 2732 2 1 2748 QDFFRBN $T=822740 769560 1 180 $X=810960 $Y=769180
X597 2519 2687 2747 2 1 2820 QDFFRBN $T=812820 799800 0 0 $X=812820 $Y=799420
X598 2499 2687 2749 2 1 2813 QDFFRBN $T=814060 819960 1 0 $X=814060 $Y=814540
X599 2833 2687 2755 2 1 2765 QDFFRBN $T=829560 830040 1 180 $X=817780 $Y=829660
X600 2773 360 2825 2 1 2850 QDFFRBN $T=819020 789720 0 0 $X=819020 $Y=789340
X601 2807 2687 2800 2 1 2841 QDFFRBN $T=823360 830040 1 0 $X=823360 $Y=824620
X602 2889 2687 2861 2 1 2817 QDFFRBN $T=840720 799800 1 180 $X=828940 $Y=799420
X603 2852 2687 2884 2 1 2843 QDFFRBN $T=830180 840120 0 0 $X=830180 $Y=839740
X604 2897 360 2825 2 1 2855 QDFFRBN $T=842580 789720 1 180 $X=830800 $Y=789340
X605 2857 2687 2884 2 1 2906 QDFFRBN $T=830800 830040 0 0 $X=830800 $Y=829660
X606 2903 2687 2749 2 1 2849 QDFFRBN $T=843820 819960 0 180 $X=832040 $Y=814540
X607 2905 360 2873 2 1 2856 QDFFRBN $T=844440 759480 1 180 $X=832660 $Y=759100
X608 2819 360 2902 2 1 2860 QDFFRBN $T=833900 779640 0 0 $X=833900 $Y=779260
X609 2874 360 2902 2 1 2921 QDFFRBN $T=835760 789720 1 0 $X=835760 $Y=784300
X610 2926 360 2873 2 1 2854 QDFFRBN $T=848160 759480 0 180 $X=836380 $Y=754060
X611 2878 2687 2800 2 1 2910 QDFFRBN $T=836380 819960 0 0 $X=836380 $Y=819580
X612 2877 2687 2861 2 1 2939 QDFFRBN $T=838860 799800 1 0 $X=838860 $Y=794380
X613 2952 360 2873 2 1 2880 QDFFRBN $T=853120 749400 1 180 $X=841340 $Y=749020
X614 2924 360 425 2 1 2888 QDFFRBN $T=853740 739320 0 180 $X=841960 $Y=733900
X615 2961 360 425 2 1 423 QDFFRBN $T=854360 719160 1 180 $X=842580 $Y=718780
X616 2962 360 425 2 1 2887 QDFFRBN $T=854360 729240 0 180 $X=842580 $Y=723820
X617 2989 2687 2861 2 1 422 QDFFRBN $T=854360 799800 1 180 $X=842580 $Y=799420
X618 2763 360 425 2 1 431 QDFFRBN $T=843200 729240 0 0 $X=843200 $Y=728860
X619 2910 2687 2914 2 1 2932 QDFFRBN $T=843820 840120 0 0 $X=843820 $Y=839740
X620 2912 2687 2914 2 1 432 QDFFRBN $T=844440 830040 0 0 $X=844440 $Y=829660
X621 2919 2687 2851 2 1 2975 QDFFRBN $T=846300 809880 0 0 $X=846300 $Y=809500
X622 2945 2687 2914 2 1 2912 QDFFRBN $T=858080 830040 0 180 $X=846300 $Y=824620
X623 2939 360 2902 2 1 3059 QDFFRBN $T=852500 789720 0 0 $X=852500 $Y=789340
X624 2973 2687 2851 2 1 3044 QDFFRBN $T=854980 819960 0 0 $X=854980 $Y=819580
X625 3016 2687 2851 2 1 2973 QDFFRBN $T=869860 809880 1 180 $X=858080 $Y=809500
X626 3013 2687 3106 2 1 3102 QDFFRBN $T=868000 799800 0 0 $X=868000 $Y=799420
X627 3129 2687 3084 2 1 3070 QDFFRBN $T=881640 819960 1 180 $X=869860 $Y=819580
X628 3031 2687 3106 2 1 3142 QDFFRBN $T=870480 799800 1 0 $X=870480 $Y=794380
X629 3080 2687 3084 2 1 460 QDFFRBN $T=871720 830040 1 0 $X=871720 $Y=824620
X630 3165 2687 3063 2 1 455 QDFFRBN $T=892800 819960 0 180 $X=881020 $Y=814540
X631 3142 2687 3106 2 1 3196 QDFFRBN $T=882260 799800 0 0 $X=882260 $Y=799420
X632 3125 2687 3106 2 1 3201 QDFFRBN $T=882260 809880 1 0 $X=882260 $Y=804460
X633 3263 2687 3221 2 1 469 QDFFRBN $T=904580 819960 0 180 $X=892800 $Y=814540
X634 3253 2687 3221 2 1 472 QDFFRBN $T=906440 809880 0 180 $X=894660 $Y=804460
X635 2567 2687 3063 2 1 3340 QDFFRBN $T=904580 819960 1 0 $X=904580 $Y=814540
X636 3385 2687 3221 2 1 495 QDFFRBN $T=928140 819960 0 180 $X=916360 $Y=814540
X637 3453 2687 3420 2 1 503 QDFFRBN $T=938060 830040 0 180 $X=926280 $Y=824620
X638 3457 2687 3425 2 1 510 QDFFRBN $T=939920 819960 0 180 $X=928140 $Y=814540
X639 2724 2687 3425 2 1 3466 QDFFRBN $T=929380 809880 1 0 $X=929380 $Y=804460
X640 2625 2687 3425 2 1 3503 QDFFRBN $T=938060 809880 0 0 $X=938060 $Y=809500
X641 3502 2687 3420 2 1 522 QDFFRBN $T=951080 830040 0 180 $X=939300 $Y=824620
X642 2719 2687 3425 2 1 3484 QDFFRBN $T=941160 819960 1 0 $X=941160 $Y=814540
X643 3568 2687 3420 2 1 536 QDFFRBN $T=966580 840120 0 180 $X=954800 $Y=834700
X644 3635 2687 3603 2 1 3617 QDFFRBN $T=981460 809880 0 180 $X=969680 $Y=804460
X645 3617 2687 3603 2 1 3642 QDFFRBN $T=971540 809880 0 0 $X=971540 $Y=809500
X646 3654 2687 3646 2 1 3635 QDFFRBN $T=993240 799800 1 180 $X=981460 $Y=799420
X647 3642 2687 3603 2 1 3656 QDFFRBN $T=982080 809880 1 0 $X=982080 $Y=804460
X648 3655 3649 3663 2 1 3666 QDFFRBN $T=992620 749400 0 0 $X=992620 $Y=749020
X649 3671 557 3661 2 1 561 QDFFRBN $T=1005640 719160 1 180 $X=993860 $Y=718780
X650 3665 557 3661 2 1 562 QDFFRBN $T=1006260 729240 0 180 $X=994480 $Y=723820
X651 3659 557 3661 2 1 3671 QDFFRBN $T=994480 729240 0 0 $X=994480 $Y=728860
X652 3657 557 3661 2 1 3665 QDFFRBN $T=994480 739320 1 0 $X=994480 $Y=733900
X653 3666 3649 3662 2 1 3657 QDFFRBN $T=1006260 749400 0 180 $X=994480 $Y=743980
X654 3667 3649 3663 2 1 3655 QDFFRBN $T=1006260 759480 0 180 $X=994480 $Y=754060
X655 3658 3649 3664 2 1 3670 QDFFRBN $T=994480 779640 0 0 $X=994480 $Y=779260
X656 3668 3649 3664 2 1 3658 QDFFRBN $T=1006260 789720 0 180 $X=994480 $Y=784300
X657 3656 2687 3646 2 1 3677 QDFFRBN $T=994480 799800 0 0 $X=994480 $Y=799420
X658 3669 3649 3646 2 1 3654 QDFFRBN $T=1006260 809880 0 180 $X=994480 $Y=804460
X659 3660 3649 3664 2 1 3667 QDFFRBN $T=995100 769560 1 0 $X=995100 $Y=764140
X660 3670 3649 3664 2 1 3660 QDFFRBN $T=1006880 769560 1 180 $X=995100 $Y=769180
X661 3673 3649 3662 2 1 3687 QDFFRBN $T=1007500 739320 0 0 $X=1007500 $Y=738940
X662 3687 3649 3663 2 1 3672 QDFFRBN $T=1019280 759480 0 180 $X=1007500 $Y=754060
X663 3672 3649 3680 2 1 3684 QDFFRBN $T=1007500 759480 0 0 $X=1007500 $Y=759100
X664 3676 3649 3646 2 1 3669 QDFFRBN $T=1019280 809880 0 180 $X=1007500 $Y=804460
X665 564 557 3661 2 1 3673 QDFFRBN $T=1019900 729240 1 180 $X=1008120 $Y=728860
X666 3683 557 3662 2 1 3659 QDFFRBN $T=1019900 739320 0 180 $X=1008120 $Y=733900
X667 3684 3649 3664 2 1 3674 QDFFRBN $T=1019900 769560 0 180 $X=1008120 $Y=764140
X668 3686 3649 3679 2 1 3668 QDFFRBN $T=1019900 789720 1 180 $X=1008120 $Y=789340
X669 3677 3649 3646 2 1 3686 QDFFRBN $T=1008120 799800 0 0 $X=1008120 $Y=799420
X670 3674 3649 3682 2 1 3685 QDFFRBN $T=1008740 779640 1 0 $X=1008740 $Y=774220
X671 3685 3649 3664 2 1 3675 QDFFRBN $T=1020520 779640 1 180 $X=1008740 $Y=779260
X672 3675 3649 3679 2 1 3691 QDFFRBN $T=1008740 789720 1 0 $X=1008740 $Y=784300
X673 3691 3649 3679 2 1 3676 QDFFRBN $T=1020520 799800 0 180 $X=1008740 $Y=794380
X674 3694 557 3678 2 1 563 QDFFRBN $T=1025480 729240 0 180 $X=1013700 $Y=723820
X675 3688 3649 3680 2 1 3698 QDFFRBN $T=1020520 759480 0 0 $X=1020520 $Y=759100
X676 3689 3649 3680 2 1 3688 QDFFRBN $T=1032920 759480 0 180 $X=1021140 $Y=754060
X677 568 3649 3662 2 1 3689 QDFFRBN $T=1033540 739320 0 180 $X=1021760 $Y=733900
X678 3692 3649 3662 2 1 3683 QDFFRBN $T=1033540 739320 1 180 $X=1021760 $Y=738940
X679 3698 3649 3682 2 1 3690 QDFFRBN $T=1033540 769560 0 180 $X=1021760 $Y=764140
X680 3704 3649 3680 2 1 3692 QDFFRBN $T=1034160 749400 0 180 $X=1022380 $Y=743980
X681 3690 3649 3682 2 1 3701 QDFFRBN $T=1022380 779640 1 0 $X=1022380 $Y=774220
X682 3695 3649 3697 2 1 3700 QDFFRBN $T=1023620 789720 1 0 $X=1023620 $Y=784300
X683 3700 3649 3679 2 1 3693 QDFFRBN $T=1035400 789720 1 180 $X=1023620 $Y=789340
X684 3693 3649 3679 2 1 3702 QDFFRBN $T=1023620 799800 1 0 $X=1023620 $Y=794380
X685 3701 3649 3696 2 1 3695 QDFFRBN $T=1036020 779640 1 180 $X=1024240 $Y=779260
X686 566 557 567 2 1 3714 QDFFRBN $T=1027960 729240 1 0 $X=1027960 $Y=723820
X687 3702 3649 3699 2 1 3703 QDFFRBN $T=1034160 799800 0 0 $X=1034160 $Y=799420
X688 3703 3649 3699 2 1 3718 QDFFRBN $T=1034780 809880 1 0 $X=1034780 $Y=804460
X689 3721 557 567 2 1 569 QDFFRBN $T=1047180 719160 1 180 $X=1035400 $Y=718780
X690 3705 557 3713 2 1 3694 QDFFRBN $T=1035400 729240 0 0 $X=1035400 $Y=728860
X691 3715 3649 3710 2 1 3705 QDFFRBN $T=1047800 739320 0 180 $X=1036020 $Y=733900
X692 3706 3649 3710 2 1 3715 QDFFRBN $T=1036640 739320 0 0 $X=1036640 $Y=738940
X693 3716 3649 3710 2 1 3704 QDFFRBN $T=1048420 749400 0 180 $X=1036640 $Y=743980
X694 3711 3649 3707 2 1 3706 QDFFRBN $T=1049040 759480 0 180 $X=1037260 $Y=754060
X695 3708 3649 3696 2 1 3723 QDFFRBN $T=1038500 769560 0 0 $X=1038500 $Y=769180
X696 3720 3649 3712 2 1 3708 QDFFRBN $T=1050280 779640 0 180 $X=1038500 $Y=774220
X697 3709 3649 3696 2 1 3720 QDFFRBN $T=1038500 779640 0 0 $X=1038500 $Y=779260
X698 3723 3649 3707 2 1 3711 QDFFRBN $T=1051520 759480 1 180 $X=1039740 $Y=759100
X699 3714 557 3713 2 1 3728 QDFFRBN $T=1042840 729240 1 0 $X=1042840 $Y=723820
X700 3717 3649 3697 2 1 3727 QDFFRBN $T=1046560 789720 0 0 $X=1046560 $Y=789340
X701 3731 3649 3697 2 1 3709 QDFFRBN $T=1058960 789720 0 180 $X=1047180 $Y=784300
X702 3729 3649 3699 2 1 3717 QDFFRBN $T=1059580 799800 0 180 $X=1047800 $Y=794380
X703 3719 3649 3699 2 1 3729 QDFFRBN $T=1047800 799800 0 0 $X=1047800 $Y=799420
X704 3718 3649 3699 2 1 3719 QDFFRBN $T=1060200 809880 0 180 $X=1048420 $Y=804460
X705 570 557 567 2 1 3721 QDFFRBN $T=1061440 719160 1 180 $X=1049660 $Y=718780
X706 3728 3649 3713 2 1 3724 QDFFRBN $T=1062060 729240 1 180 $X=1050280 $Y=728860
X707 3724 3649 3713 2 1 3725 QDFFRBN $T=1050900 739320 1 0 $X=1050900 $Y=733900
X708 3725 3649 3722 2 1 3737 QDFFRBN $T=1050900 739320 0 0 $X=1050900 $Y=738940
X709 3733 3649 3722 2 1 3716 QDFFRBN $T=1062680 749400 1 180 $X=1050900 $Y=749020
X710 3726 3649 3722 2 1 3733 QDFFRBN $T=1050900 759480 1 0 $X=1050900 $Y=754060
X711 3732 3649 3712 2 1 3726 QDFFRBN $T=1063300 769560 0 180 $X=1051520 $Y=764140
X712 3727 3649 3730 2 1 3732 QDFFRBN $T=1051520 769560 0 0 $X=1051520 $Y=769180
X713 3741 3649 3697 2 1 3731 QDFFRBN $T=1072600 789720 0 180 $X=1060820 $Y=784300
X714 3737 3649 3722 2 1 3742 QDFFRBN $T=1064540 739320 0 0 $X=1064540 $Y=738940
X715 3742 3649 3722 2 1 3734 QDFFRBN $T=1076940 749400 0 180 $X=1065160 $Y=743980
X716 3734 3649 3722 2 1 3735 QDFFRBN $T=1076940 749400 1 180 $X=1065160 $Y=749020
X717 3735 3649 3730 2 1 3738 QDFFRBN $T=1065160 759480 1 0 $X=1065160 $Y=754060
X718 3738 3649 3730 2 1 3744 QDFFRBN $T=1065160 759480 0 0 $X=1065160 $Y=759100
X719 3739 3649 3730 2 1 3743 QDFFRBN $T=1065160 769560 0 0 $X=1065160 $Y=769180
X720 3743 3649 3730 2 1 3736 QDFFRBN $T=1076940 779640 1 180 $X=1065160 $Y=779260
X721 3744 3649 3730 2 1 3739 QDFFRBN $T=1077560 769560 0 180 $X=1065780 $Y=764140
X722 3736 3649 3740 2 1 3745 QDFFRBN $T=1066400 799800 1 0 $X=1066400 $Y=794380
X723 3745 3649 3740 2 1 3741 QDFFRBN $T=1078800 789720 1 180 $X=1067020 $Y=789340
X724 599 2 592 1 INV1S $T=311240 759480 0 180 $X=310000 $Y=754060
X725 604 2 601 1 INV1S $T=315580 739320 0 180 $X=314340 $Y=733900
X726 611 2 598 1 INV1S $T=319300 789720 1 180 $X=318060 $Y=789340
X727 603 2 612 1 INV1S $T=318680 749400 0 0 $X=318680 $Y=749020
X728 624 2 616 1 INV1S $T=322400 739320 1 180 $X=321160 $Y=738940
X729 645 2 634 1 INV1S $T=327980 749400 0 180 $X=326740 $Y=743980
X730 626 2 639 1 INV1S $T=328600 799800 1 180 $X=327360 $Y=799420
X731 595 2 614 1 INV1S $T=328600 809880 0 180 $X=327360 $Y=804460
X732 653 2 595 1 INV1S $T=329840 809880 0 180 $X=328600 $Y=804460
X733 636 2 648 1 INV1S $T=332320 739320 1 180 $X=331080 $Y=738940
X734 643 2 660 1 INV1S $T=333560 779640 1 180 $X=332320 $Y=779260
X735 635 2 661 1 INV1S $T=334180 729240 1 180 $X=332940 $Y=728860
X736 679 2 680 1 INV1S $T=337280 809880 0 180 $X=336040 $Y=804460
X737 686 2 673 1 INV1S $T=337900 759480 1 180 $X=336660 $Y=759100
X738 687 2 686 1 INV1S $T=339140 759480 1 180 $X=337900 $Y=759100
X739 693 2 699 1 INV1S $T=339140 749400 0 0 $X=339140 $Y=749020
X740 696 2 668 1 INV1S $T=340380 759480 1 180 $X=339140 $Y=759100
X741 695 2 696 1 INV1S $T=341620 759480 1 180 $X=340380 $Y=759100
X742 713 2 689 1 INV1S $T=342860 799800 0 180 $X=341620 $Y=794380
X743 719 2 713 1 INV1S $T=345960 799800 1 0 $X=345960 $Y=794380
X744 749 2 722 1 INV1S $T=349680 769560 0 180 $X=348440 $Y=764140
X745 732 2 710 1 INV1S $T=350920 749400 1 180 $X=349680 $Y=749020
X746 745 2 751 1 INV1S $T=355260 779640 0 0 $X=355260 $Y=779260
X747 744 2 755 1 INV1S $T=357740 759480 0 0 $X=357740 $Y=759100
X748 22 2 23 1 INV1S $T=360220 719160 0 0 $X=360220 $Y=718780
X749 763 2 721 1 INV1S $T=362700 729240 1 180 $X=361460 $Y=728860
X750 767 2 757 1 INV1S $T=363320 739320 0 180 $X=362080 $Y=733900
X751 741 2 771 1 INV1S $T=362080 890520 0 0 $X=362080 $Y=890140
X752 783 2 774 1 INV1S $T=366420 769560 0 180 $X=365180 $Y=764140
X753 795 2 778 1 INV1S $T=367040 799800 1 180 $X=365800 $Y=799420
X754 784 2 793 1 INV1S $T=369520 789720 0 180 $X=368280 $Y=784300
X755 750 2 807 1 INV1S $T=369520 880440 0 0 $X=369520 $Y=880060
X756 812 2 800 1 INV1S $T=371380 779640 1 180 $X=370140 $Y=779260
X757 817 2 786 1 INV1S $T=371380 809880 0 180 $X=370140 $Y=804460
X758 815 2 811 1 INV1S $T=372000 749400 0 180 $X=370760 $Y=743980
X759 816 2 799 1 INV1S $T=372000 759480 1 180 $X=370760 $Y=759100
X760 826 2 819 1 INV1S $T=376960 739320 0 180 $X=375720 $Y=733900
X761 825 2 818 1 INV1S $T=377580 729240 0 180 $X=376340 $Y=723820
X762 832 2 821 1 INV1S $T=377580 789720 1 180 $X=376340 $Y=789340
X763 830 2 838 1 INV1S $T=377580 759480 1 0 $X=377580 $Y=754060
X764 835 2 836 1 INV1S $T=377580 880440 1 0 $X=377580 $Y=875020
X765 838 2 828 1 INV1S $T=379440 769560 0 180 $X=378200 $Y=764140
X766 838 2 775 1 INV1S $T=378820 779640 1 0 $X=378820 $Y=774220
X767 844 2 849 1 INV1S $T=379440 729240 0 0 $X=379440 $Y=728860
X768 39 2 35 1 INV1S $T=380060 900600 1 0 $X=380060 $Y=895180
X769 863 2 860 1 INV1S $T=383160 759480 1 180 $X=381920 $Y=759100
X770 846 2 840 1 INV1S $T=383160 769560 0 180 $X=381920 $Y=764140
X771 859 2 823 1 INV1S $T=381920 890520 0 0 $X=381920 $Y=890140
X772 861 2 877 1 INV1S $T=383780 860280 0 0 $X=383780 $Y=859900
X773 870 2 852 1 INV1S $T=384400 749400 1 0 $X=384400 $Y=743980
X774 879 2 885 1 INV1S $T=385020 850200 0 0 $X=385020 $Y=849820
X775 875 2 881 1 INV1S $T=386880 729240 1 180 $X=385640 $Y=728860
X776 887 2 876 1 INV1S $T=386260 870360 1 0 $X=386260 $Y=864940
X777 854 2 903 1 INV1S $T=386880 779640 0 0 $X=386880 $Y=779260
X778 872 2 867 1 INV1S $T=387500 840120 1 0 $X=387500 $Y=834700
X779 901 2 898 1 INV1S $T=389360 789720 1 180 $X=388120 $Y=789340
X780 904 2 871 1 INV1S $T=389980 759480 1 180 $X=388740 $Y=759100
X781 891 2 910 1 INV1S $T=389980 719160 0 0 $X=389980 $Y=718780
X782 909 2 848 1 INV1S $T=391840 890520 0 180 $X=390600 $Y=885100
X783 857 2 908 1 INV1S $T=391220 779640 1 0 $X=391220 $Y=774220
X784 949 2 43 1 INV1S $T=393700 900600 0 180 $X=392460 $Y=895180
X785 928 2 916 1 INV1S $T=398040 840120 0 0 $X=398040 $Y=839740
X786 944 2 932 1 INV1S $T=399280 860280 0 180 $X=398040 $Y=854860
X787 938 2 880 1 INV1S $T=398660 880440 0 0 $X=398660 $Y=880060
X788 45 2 953 1 INV1S $T=399280 870360 0 0 $X=399280 $Y=869980
X789 961 2 946 1 INV1S $T=402380 769560 1 180 $X=401140 $Y=769180
X790 54 2 954 1 INV1S $T=403000 900600 0 180 $X=401760 $Y=895180
X791 976 2 961 1 INV1S $T=404240 769560 1 180 $X=403000 $Y=769180
X792 950 2 963 1 INV1S $T=404860 759480 1 180 $X=403620 $Y=759100
X793 924 2 969 1 INV1S $T=403620 819960 0 0 $X=403620 $Y=819580
X794 980 2 958 1 INV1S $T=406720 729240 1 180 $X=405480 $Y=728860
X795 988 2 900 1 INV1S $T=407340 880440 0 180 $X=406100 $Y=875020
X796 912 2 985 1 INV1S $T=406720 749400 0 0 $X=406720 $Y=749020
X797 1000 2 951 1 INV1S $T=407960 840120 0 180 $X=406720 $Y=834700
X798 941 2 993 1 INV1S $T=407960 769560 1 0 $X=407960 $Y=764140
X799 920 2 999 1 INV1S $T=407960 799800 0 0 $X=407960 $Y=799420
X800 1009 2 966 1 INV1S $T=410440 880440 0 180 $X=409200 $Y=875020
X801 1004 2 1010 1 INV1S $T=410440 819960 1 0 $X=410440 $Y=814540
X802 1001 2 986 1 INV1S $T=413540 739320 0 180 $X=412300 $Y=733900
X803 998 2 1020 1 INV1S $T=412920 789720 1 0 $X=412920 $Y=784300
X804 1023 2 1038 1 INV1S $T=413540 850200 0 0 $X=413540 $Y=849820
X805 967 2 1018 1 INV1S $T=415400 769560 0 180 $X=414160 $Y=764140
X806 1024 2 990 1 INV1S $T=414160 860280 0 0 $X=414160 $Y=859900
X807 973 2 62 1 INV1S $T=417260 739320 1 180 $X=416020 $Y=738940
X808 1026 2 65 1 INV1S $T=417260 900600 1 0 $X=417260 $Y=895180
X809 1036 2 1037 1 INV1S $T=418500 809880 0 0 $X=418500 $Y=809500
X810 1043 2 1042 1 INV1S $T=419740 890520 0 0 $X=419740 $Y=890140
X811 1046 2 1031 1 INV1S $T=420360 779640 1 0 $X=420360 $Y=774220
X812 1019 2 1047 1 INV1S $T=420360 840120 1 0 $X=420360 $Y=834700
X813 1051 2 1005 1 INV1S $T=422220 819960 1 180 $X=420980 $Y=819580
X814 1035 2 1049 1 INV1S $T=423460 739320 1 0 $X=423460 $Y=733900
X815 1068 2 1053 1 INV1S $T=425940 860280 1 180 $X=424700 $Y=859900
X816 1069 2 1030 1 INV1S $T=425940 880440 0 180 $X=424700 $Y=875020
X817 834 2 1073 1 INV1S $T=427180 789720 1 0 $X=427180 $Y=784300
X818 72 2 1088 1 INV1S $T=428420 729240 1 0 $X=428420 $Y=723820
X819 1054 2 1087 1 INV1S $T=430900 809880 1 0 $X=430900 $Y=804460
X820 1066 2 1080 1 INV1S $T=430900 850200 0 0 $X=430900 $Y=849820
X821 1086 2 1093 1 INV1S $T=431520 759480 0 0 $X=431520 $Y=759100
X822 1105 2 1063 1 INV1S $T=434620 830040 1 180 $X=433380 $Y=829660
X823 1050 2 1109 1 INV1S $T=434620 739320 0 0 $X=434620 $Y=738940
X824 1102 2 74 1 INV1S $T=434620 890520 1 0 $X=434620 $Y=885100
X825 1100 2 77 1 INV1S $T=435860 900600 0 180 $X=434620 $Y=895180
X826 1052 2 1108 1 INV1S $T=435240 759480 1 0 $X=435240 $Y=754060
X827 1081 2 1123 1 INV1S $T=437100 860280 0 0 $X=437100 $Y=859900
X828 1072 2 1099 1 INV1S $T=438960 759480 0 180 $X=437720 $Y=754060
X829 1127 2 1071 1 INV1S $T=442680 749400 1 180 $X=441440 $Y=749020
X830 1132 2 1127 1 INV1S $T=443300 749400 0 180 $X=442060 $Y=743980
X831 1150 2 1112 1 INV1S $T=445160 840120 1 180 $X=443920 $Y=839740
X832 1140 2 1116 1 INV1S $T=443920 880440 0 0 $X=443920 $Y=880060
X833 1121 2 1143 1 INV1S $T=444540 860280 1 0 $X=444540 $Y=854860
X834 1139 2 1115 1 INV1S $T=444540 870360 0 0 $X=444540 $Y=869980
X835 1147 2 1091 1 INV1S $T=447020 890520 0 180 $X=445780 $Y=885100
X836 1146 2 92 1 INV1S $T=446400 719160 0 0 $X=446400 $Y=718780
X837 1125 2 1148 1 INV1S $T=446400 729240 0 0 $X=446400 $Y=728860
X838 1155 2 1134 1 INV1S $T=448880 799800 1 180 $X=447640 $Y=799420
X839 1178 2 1089 1 INV1S $T=448880 819960 1 180 $X=447640 $Y=819580
X840 1142 2 1149 1 INV1S $T=448880 799800 0 0 $X=448880 $Y=799420
X841 1159 2 1152 1 INV1S $T=450120 880440 1 180 $X=448880 $Y=880060
X842 1158 2 96 1 INV1S $T=448880 890520 0 0 $X=448880 $Y=890140
X843 1168 2 1124 1 INV1S $T=451980 789720 0 0 $X=451980 $Y=789340
X844 1173 2 1162 1 INV1S $T=453220 860280 0 180 $X=451980 $Y=854860
X845 1175 2 1151 1 INV1S $T=453220 870360 0 180 $X=451980 $Y=864940
X846 1169 2 1174 1 INV1S $T=453220 840120 1 0 $X=453220 $Y=834700
X847 1182 2 1145 1 INV1S $T=455700 789720 0 180 $X=454460 $Y=784300
X848 1179 2 1184 1 INV1S $T=455080 779640 0 0 $X=455080 $Y=779260
X849 1156 2 1185 1 INV1S $T=456320 819960 1 0 $X=456320 $Y=814540
X850 1180 2 1195 1 INV1S $T=458180 850200 1 0 $X=458180 $Y=844780
X851 1202 2 1113 1 INV1S $T=461280 799800 1 180 $X=460040 $Y=799420
X852 1207 2 1177 1 INV1S $T=462520 880440 1 180 $X=461280 $Y=880060
X853 1190 2 1210 1 INV1S $T=462520 799800 0 0 $X=462520 $Y=799420
X854 1181 2 1215 1 INV1S $T=463140 870360 1 0 $X=463140 $Y=864940
X855 1186 2 1203 1 INV1S $T=463760 830040 0 0 $X=463760 $Y=829660
X856 1231 2 1216 1 INV1S $T=467480 819960 0 180 $X=466240 $Y=814540
X857 1223 2 1211 1 INV1S $T=469340 769560 0 0 $X=469340 $Y=769180
X858 1253 2 1229 1 INV1S $T=471820 830040 1 180 $X=470580 $Y=829660
X859 1224 2 1209 1 INV1S $T=472440 729240 1 180 $X=471200 $Y=728860
X860 1244 2 103 1 INV1S $T=472440 890520 1 180 $X=471200 $Y=890140
X861 1247 2 1246 1 INV1S $T=472440 850200 0 0 $X=472440 $Y=849820
X862 1249 2 1228 1 INV1S $T=474300 890520 1 180 $X=473060 $Y=890140
X863 1261 2 1258 1 INV1S $T=476160 759480 1 0 $X=476160 $Y=754060
X864 1268 2 1240 1 INV1S $T=477400 860280 1 180 $X=476160 $Y=859900
X865 1283 2 1271 1 INV1S $T=479260 840120 1 180 $X=478020 $Y=839740
X866 1273 2 1272 1 INV1S $T=478020 880440 1 0 $X=478020 $Y=875020
X867 1267 2 1270 1 INV1S $T=478640 759480 1 0 $X=478640 $Y=754060
X868 1294 2 1274 1 INV1S $T=481740 850200 0 180 $X=480500 $Y=844780
X869 1295 2 1276 1 INV1S $T=482980 729240 1 180 $X=481740 $Y=728860
X870 1302 2 1254 1 INV1S $T=482980 819960 0 180 $X=481740 $Y=814540
X871 1289 2 1260 1 INV1S $T=482980 789720 0 0 $X=482980 $Y=789340
X872 1310 2 1307 1 INV1S $T=484840 890520 0 0 $X=484840 $Y=890140
X873 127 2 1265 1 INV1S $T=487320 739320 1 180 $X=486080 $Y=738940
X874 1311 2 1305 1 INV1S $T=486700 799800 1 0 $X=486700 $Y=794380
X875 1301 2 1236 1 INV1S $T=487940 819960 0 180 $X=486700 $Y=814540
X876 1323 2 1280 1 INV1S $T=487940 830040 1 180 $X=486700 $Y=829660
X877 1306 2 1309 1 INV1S $T=488560 830040 1 0 $X=488560 $Y=824620
X878 1324 2 1288 1 INV1S $T=489180 779640 0 0 $X=489180 $Y=779260
X879 129 2 1281 1 INV1S $T=491040 739320 1 180 $X=489800 $Y=738940
X880 1342 2 1313 1 INV1S $T=491660 769560 1 180 $X=490420 $Y=769180
X881 1340 2 1285 1 INV1S $T=491660 860280 1 180 $X=490420 $Y=859900
X882 1296 2 1331 1 INV1S $T=490420 880440 1 0 $X=490420 $Y=875020
X883 1333 2 1297 1 INV1S $T=492900 739320 0 180 $X=491660 $Y=733900
X884 134 2 1279 1 INV1S $T=493520 739320 1 180 $X=492280 $Y=738940
X885 1348 2 1316 1 INV1S $T=494760 860280 1 180 $X=493520 $Y=859900
X886 1341 2 1327 1 INV1S $T=493520 880440 0 0 $X=493520 $Y=880060
X887 136 2 126 1 INV1S $T=495380 719160 1 180 $X=494140 $Y=718780
X888 1366 2 1278 1 INV1S $T=496000 739320 1 180 $X=494760 $Y=738940
X889 1362 2 1318 1 INV1S $T=496620 729240 1 180 $X=495380 $Y=728860
X890 1357 2 1349 1 INV1S $T=496620 850200 1 180 $X=495380 $Y=849820
X891 137 2 138 1 INV1S $T=496000 719160 0 0 $X=496000 $Y=718780
X892 1358 2 1130 1 INV1S $T=497240 890520 0 180 $X=496000 $Y=885100
X893 1361 2 1351 1 INV1S $T=499100 890520 1 180 $X=497860 $Y=890140
X894 1370 2 1356 1 INV1S $T=500340 840120 0 180 $X=499100 $Y=834700
X895 1380 2 1359 1 INV1S $T=500960 769560 1 180 $X=499720 $Y=769180
X896 1376 2 1300 1 INV1S $T=502200 779640 0 180 $X=500960 $Y=774220
X897 1354 2 1379 1 INV1S $T=501580 860280 0 0 $X=501580 $Y=859900
X898 1375 2 1343 1 INV1S $T=502200 759480 1 0 $X=502200 $Y=754060
X899 1371 2 1335 1 INV1S $T=502200 799800 0 0 $X=502200 $Y=799420
X900 1372 2 143 1 INV1S $T=502200 900600 1 0 $X=502200 $Y=895180
X901 1389 2 1329 1 INV1S $T=504060 799800 0 180 $X=502820 $Y=794380
X902 1392 2 1384 1 INV1S $T=504680 809880 0 180 $X=503440 $Y=804460
X903 1377 2 1385 1 INV1S $T=504060 819960 1 0 $X=504060 $Y=814540
X904 1383 2 1314 1 INV1S $T=505920 789720 0 0 $X=505920 $Y=789340
X905 1399 2 1365 1 INV1S $T=507160 870360 0 180 $X=505920 $Y=864940
X906 1398 2 1388 1 INV1S $T=505920 890520 1 0 $X=505920 $Y=885100
X907 1403 2 1364 1 INV1S $T=507780 840120 0 180 $X=506540 $Y=834700
X908 1397 2 1421 1 INV1S $T=507780 880440 1 0 $X=507780 $Y=875020
X909 1378 2 1409 1 INV1S $T=508400 830040 1 0 $X=508400 $Y=824620
X910 1428 2 1393 1 INV1S $T=512740 729240 1 180 $X=511500 $Y=728860
X911 152 2 1406 1 INV1S $T=512740 900600 0 180 $X=511500 $Y=895180
X912 1427 2 1401 1 INV1S $T=513360 779640 0 180 $X=512120 $Y=774220
X913 1415 2 1417 1 INV1S $T=512120 809880 1 0 $X=512120 $Y=804460
X914 1434 2 1426 1 INV1S $T=514600 769560 0 180 $X=513360 $Y=764140
X915 1358 2 146 1 INV1S $T=513980 739320 0 0 $X=513980 $Y=738940
X916 1431 2 1412 1 INV1S $T=515840 749400 0 180 $X=514600 $Y=743980
X917 1408 2 155 1 INV1S $T=515220 870360 0 0 $X=515220 $Y=869980
X918 1443 2 1416 1 INV1S $T=516460 890520 1 0 $X=516460 $Y=885100
X919 1453 2 1438 1 INV1S $T=518320 759480 1 180 $X=517080 $Y=759100
X920 1449 2 1423 1 INV1S $T=518320 840120 0 0 $X=518320 $Y=839740
X921 1451 2 1418 1 INV1S $T=520180 880440 1 180 $X=518940 $Y=880060
X922 1454 2 1432 1 INV1S $T=520180 850200 0 0 $X=520180 $Y=849820
X923 1466 2 1448 1 INV1S $T=522040 860280 1 180 $X=520800 $Y=859900
X924 1469 2 1437 1 INV1S $T=522660 729240 1 180 $X=521420 $Y=728860
X925 1429 2 1463 1 INV1S $T=521420 799800 1 0 $X=521420 $Y=794380
X926 162 2 1452 1 INV1S $T=523900 900600 0 180 $X=522660 $Y=895180
X927 1473 2 1464 1 INV1S $T=523900 830040 0 0 $X=523900 $Y=829660
X928 1457 2 1336 1 INV1S $T=525760 769560 0 180 $X=524520 $Y=764140
X929 1460 2 1489 1 INV1S $T=525760 850200 1 0 $X=525760 $Y=844780
X930 1481 2 1485 1 INV1S $T=526380 789720 1 0 $X=526380 $Y=784300
X931 1509 2 1476 1 INV1S $T=528860 769560 0 180 $X=527620 $Y=764140
X932 1439 2 1479 1 INV1S $T=528240 819960 0 0 $X=528240 $Y=819580
X933 1487 2 1413 1 INV1S $T=528860 779640 0 0 $X=528860 $Y=779260
X934 1500 2 1450 1 INV1S $T=530100 880440 1 180 $X=528860 $Y=880060
X935 1513 2 1494 1 INV1S $T=531960 860280 1 180 $X=530720 $Y=859900
X936 1492 2 1503 1 INV1S $T=532580 799800 0 180 $X=531340 $Y=794380
X937 1493 2 1520 1 INV1S $T=531960 819960 1 0 $X=531960 $Y=814540
X938 1515 2 1499 1 INV1S $T=533200 830040 0 180 $X=531960 $Y=824620
X939 1518 2 1502 1 INV1S $T=534440 890520 1 180 $X=533200 $Y=890140
X940 1517 2 1498 1 INV1S $T=533820 840120 1 0 $X=533820 $Y=834700
X941 1507 2 167 1 INV1S $T=535060 729240 1 0 $X=535060 $Y=723820
X942 1506 2 169 1 INV1S $T=535060 880440 1 0 $X=535060 $Y=875020
X943 1525 2 1514 1 INV1S $T=536300 850200 0 0 $X=536300 $Y=849820
X944 1531 2 1488 1 INV1S $T=537540 880440 1 0 $X=537540 $Y=875020
X945 1538 2 1526 1 INV1S $T=539400 789720 1 180 $X=538160 $Y=789340
X946 1548 2 1470 1 INV1S $T=540020 729240 0 180 $X=538780 $Y=723820
X947 1532 2 1455 1 INV1S $T=538780 749400 1 0 $X=538780 $Y=743980
X948 1542 2 1510 1 INV1S $T=540020 779640 1 180 $X=538780 $Y=779260
X949 1533 2 1480 1 INV1S $T=538780 890520 1 0 $X=538780 $Y=885100
X950 1522 2 1550 1 INV1S $T=540020 819960 0 0 $X=540020 $Y=819580
X951 1555 2 1530 1 INV1S $T=541880 860280 1 180 $X=540640 $Y=859900
X952 1557 2 1535 1 INV1S $T=542500 749400 0 180 $X=541260 $Y=743980
X953 1534 2 1536 1 INV1S $T=543120 779640 1 0 $X=543120 $Y=774220
X954 1568 2 1546 1 INV1S $T=544980 840120 0 180 $X=543740 $Y=834700
X955 1559 2 1528 1 INV1S $T=544360 759480 1 0 $X=544360 $Y=754060
X956 1573 2 1539 1 INV1S $T=546220 840120 1 180 $X=544980 $Y=839740
X957 1581 2 1584 1 INV1S $T=547460 759480 0 0 $X=547460 $Y=759100
X958 1592 2 1566 1 INV1S $T=548700 789720 1 180 $X=547460 $Y=789340
X959 174 2 1547 1 INV1S $T=548700 900600 0 180 $X=547460 $Y=895180
X960 1588 2 1574 1 INV1S $T=549320 890520 0 180 $X=548080 $Y=885100
X961 1578 2 1582 1 INV1S $T=548700 850200 0 0 $X=548700 $Y=849820
X962 1614 2 1497 1 INV1S $T=551800 830040 0 180 $X=550560 $Y=824620
X963 1590 2 173 1 INV1S $T=551180 729240 1 0 $X=551180 $Y=723820
X964 1601 2 1585 1 INV1S $T=552420 860280 1 180 $X=551180 $Y=859900
X965 1591 2 1543 1 INV1S $T=551800 779640 1 0 $X=551800 $Y=774220
X966 1607 2 1593 1 INV1S $T=554280 880440 0 180 $X=553040 $Y=875020
X967 1608 2 1565 1 INV1S $T=555520 729240 0 180 $X=554280 $Y=723820
X968 1625 2 1549 1 INV1S $T=555520 789720 1 180 $X=554280 $Y=789340
X969 1603 2 1577 1 INV1S $T=555520 749400 0 0 $X=555520 $Y=749020
X970 1605 2 1567 1 INV1S $T=555520 809880 1 0 $X=555520 $Y=804460
X971 1612 2 1529 1 INV1S $T=556760 779640 0 0 $X=556760 $Y=779260
X972 135 2 176 1 INV1S $T=557380 729240 1 0 $X=557380 $Y=723820
X973 1616 2 1586 1 INV1S $T=557380 799800 1 0 $X=557380 $Y=794380
X974 1611 2 1587 1 INV1S $T=558000 739320 0 0 $X=558000 $Y=738940
X975 1631 2 1627 1 INV1S $T=558620 759480 1 0 $X=558620 $Y=754060
X976 1634 2 1639 1 INV1S $T=559240 789720 0 0 $X=559240 $Y=789340
X977 1645 2 1610 1 INV1S $T=561100 850200 0 180 $X=559860 $Y=844780
X978 1630 2 1628 1 INV1S $T=560480 860280 0 0 $X=560480 $Y=859900
X979 1655 2 1638 1 INV1S $T=564820 840120 1 180 $X=563580 $Y=839740
X980 1670 2 1641 1 INV1S $T=568540 729240 0 180 $X=567300 $Y=723820
X981 1677 2 1657 1 INV1S $T=569160 860280 1 180 $X=567920 $Y=859900
X982 1678 2 1637 1 INV1S $T=569160 880440 0 180 $X=567920 $Y=875020
X983 1663 2 1604 1 INV1S $T=567920 890520 1 0 $X=567920 $Y=885100
X984 1665 2 1640 1 INV1S $T=568540 729240 0 0 $X=568540 $Y=728860
X985 1683 2 1654 1 INV1S $T=569780 769560 0 180 $X=568540 $Y=764140
X986 1676 2 1651 1 INV1S $T=569780 830040 1 180 $X=568540 $Y=829660
X987 1681 2 1644 1 INV1S $T=570400 900600 0 180 $X=569160 $Y=895180
X988 1687 2 1656 1 INV1S $T=571020 739320 1 180 $X=569780 $Y=738940
X989 1693 2 1662 1 INV1S $T=571640 799800 0 180 $X=570400 $Y=794380
X990 1675 2 1594 1 INV1S $T=570400 809880 1 0 $X=570400 $Y=804460
X991 1672 2 1598 1 INV1S $T=572260 809880 1 180 $X=571020 $Y=809500
X992 1700 2 1624 1 INV1S $T=574120 779640 0 0 $X=574120 $Y=779260
X993 1706 2 1692 1 INV1S $T=575360 870360 1 180 $X=574120 $Y=869980
X994 1695 2 1679 1 INV1S $T=575360 739320 1 0 $X=575360 $Y=733900
X995 1716 2 1696 1 INV1S $T=577220 830040 0 180 $X=575980 $Y=824620
X996 1720 2 1684 1 INV1S $T=578460 840120 1 180 $X=577220 $Y=839740
X997 1724 2 1664 1 INV1S $T=578460 860280 0 180 $X=577220 $Y=854860
X998 1725 2 1658 1 INV1S $T=579700 749400 0 180 $X=578460 $Y=743980
X999 1685 2 1721 1 INV1S $T=578460 890520 1 0 $X=578460 $Y=885100
X1000 1741 2 1708 1 INV1S $T=580940 749400 1 180 $X=579700 $Y=749020
X1001 1739 2 1712 1 INV1S $T=582800 779640 0 180 $X=581560 $Y=774220
X1002 1742 2 1702 1 INV1S $T=583420 870360 0 0 $X=583420 $Y=869980
X1003 1746 2 1729 1 INV1S $T=584040 779640 0 0 $X=584040 $Y=779260
X1004 1771 2 1709 1 INV1S $T=585280 840120 1 180 $X=584040 $Y=839740
X1005 1756 2 1731 1 INV1S $T=586520 830040 0 180 $X=585280 $Y=824620
X1006 1758 2 1738 1 INV1S $T=587760 729240 1 180 $X=586520 $Y=728860
X1007 1753 2 1713 1 INV1S $T=586520 799800 1 0 $X=586520 $Y=794380
X1008 1757 2 1732 1 INV1S $T=587140 870360 0 0 $X=587140 $Y=869980
X1009 1764 2 1691 1 INV1S $T=588380 769560 1 0 $X=588380 $Y=764140
X1010 1770 2 1747 1 INV1S $T=590240 799800 0 180 $X=589000 $Y=794380
X1011 1774 2 1755 1 INV1S $T=590860 880440 0 0 $X=590860 $Y=880060
X1012 1768 2 1773 1 INV1S $T=591480 860280 0 0 $X=591480 $Y=859900
X1013 1777 2 1719 1 INV1S $T=593960 809880 0 0 $X=593960 $Y=809500
X1014 1785 2 1788 1 INV1S $T=594580 789720 0 0 $X=594580 $Y=789340
X1015 1782 2 1779 1 INV1S $T=594580 830040 1 0 $X=594580 $Y=824620
X1016 1786 2 1735 1 INV1S $T=597680 840120 0 180 $X=596440 $Y=834700
X1017 1805 2 1765 1 INV1S $T=598920 779640 0 180 $X=597680 $Y=774220
X1018 1800 2 1754 1 INV1S $T=598920 819960 1 180 $X=597680 $Y=819580
X1019 1763 2 1803 1 INV1S $T=598300 850200 1 0 $X=598300 $Y=844780
X1020 1813 2 1767 1 INV1S $T=600160 749400 1 180 $X=598920 $Y=749020
X1021 1815 2 1789 1 INV1S $T=600160 870360 1 180 $X=598920 $Y=869980
X1022 1809 2 1804 1 INV1S $T=600160 880440 1 180 $X=598920 $Y=880060
X1023 1806 2 191 1 INV1S $T=601400 719160 1 180 $X=600160 $Y=718780
X1024 1816 2 1761 1 INV1S $T=601400 779640 0 180 $X=600160 $Y=774220
X1025 1821 2 1766 1 INV1S $T=602020 749400 0 180 $X=600780 $Y=743980
X1026 1807 2 1819 1 INV1S $T=601400 759480 0 0 $X=601400 $Y=759100
X1027 1829 2 1808 1 INV1S $T=605120 789720 1 180 $X=603880 $Y=789340
X1028 1835 2 1795 1 INV1S $T=605120 809880 1 180 $X=603880 $Y=809500
X1029 1843 2 1823 1 INV1S $T=606360 890520 0 180 $X=605120 $Y=885100
X1030 1849 2 1824 1 INV1S $T=607600 779640 0 180 $X=606360 $Y=774220
X1031 1844 2 1841 1 INV1S $T=607600 809880 1 180 $X=606360 $Y=809500
X1032 1845 2 1812 1 INV1S $T=607600 830040 0 180 $X=606360 $Y=824620
X1033 206 2 202 1 INV1S $T=608840 719160 1 180 $X=607600 $Y=718780
X1034 1854 2 1797 1 INV1S $T=609460 749400 1 180 $X=608220 $Y=749020
X1035 1850 2 1836 1 INV1S $T=608220 840120 1 0 $X=608220 $Y=834700
X1036 1820 2 1855 1 INV1S $T=608840 799800 1 0 $X=608840 $Y=794380
X1037 1860 2 1830 1 INV1S $T=610080 850200 0 180 $X=608840 $Y=844780
X1038 1861 2 1831 1 INV1S $T=610080 870360 0 180 $X=608840 $Y=864940
X1039 1838 2 1873 1 INV1S $T=611320 799800 1 0 $X=611320 $Y=794380
X1040 1866 2 1801 1 INV1S $T=613180 860280 0 0 $X=613180 $Y=859900
X1041 209 2 1653 1 INV1S $T=615040 739320 0 180 $X=613800 $Y=733900
X1042 1877 2 208 1 INV1S $T=616280 729240 1 180 $X=615040 $Y=728860
X1043 1875 2 1847 1 INV1S $T=616280 749400 0 180 $X=615040 $Y=743980
X1044 1882 2 1794 1 INV1S $T=616280 739320 0 0 $X=616280 $Y=738940
X1045 1896 2 1880 1 INV1S $T=617520 860280 1 180 $X=616280 $Y=859900
X1046 1891 2 1885 1 INV1S $T=618760 749400 1 180 $X=617520 $Y=749020
X1047 1888 2 1895 1 INV1S $T=617520 789720 0 0 $X=617520 $Y=789340
X1048 1890 2 1832 1 INV1S $T=618760 880440 1 180 $X=617520 $Y=880060
X1049 1848 2 1892 1 INV1S $T=618140 809880 1 0 $X=618140 $Y=804460
X1050 1900 2 1879 1 INV1S $T=620000 850200 0 180 $X=618760 $Y=844780
X1051 1893 2 1897 1 INV1S $T=618760 880440 0 0 $X=618760 $Y=880060
X1052 1905 2 1865 1 INV1S $T=620620 900600 0 180 $X=619380 $Y=895180
X1053 1908 2 1862 1 INV1S $T=621240 769560 0 180 $X=620000 $Y=764140
X1054 1902 2 1876 1 INV1S $T=621240 840120 0 180 $X=620000 $Y=834700
X1055 1924 2 1878 1 INV1S $T=622480 819960 1 180 $X=621240 $Y=819580
X1056 1903 2 1870 1 INV1S $T=621860 830040 0 0 $X=621860 $Y=829660
X1057 1898 2 1913 1 INV1S $T=622480 779640 1 0 $X=622480 $Y=774220
X1058 217 2 216 1 INV1S $T=623720 900600 0 180 $X=622480 $Y=895180
X1059 199 2 1833 1 INV1S $T=623100 759480 0 0 $X=623100 $Y=759100
X1060 1916 2 214 1 INV1S $T=623720 729240 1 0 $X=623720 $Y=723820
X1061 1935 2 212 1 INV1S $T=627440 739320 0 180 $X=626200 $Y=733900
X1062 1936 2 1923 1 INV1S $T=627440 809880 0 180 $X=626200 $Y=804460
X1063 1919 2 1846 1 INV1S $T=626820 860280 1 0 $X=626820 $Y=854860
X1064 1927 2 1950 1 INV1S $T=631160 819960 0 0 $X=631160 $Y=819580
X1065 1934 2 1945 1 INV1S $T=631780 799800 0 0 $X=631780 $Y=799420
X1066 1960 2 1928 1 INV1S $T=633020 890520 0 180 $X=631780 $Y=885100
X1067 1963 2 1933 1 INV1S $T=633640 769560 1 180 $X=632400 $Y=769180
X1068 225 2 218 1 INV1S $T=633640 900600 0 180 $X=632400 $Y=895180
X1069 1967 2 1899 1 INV1S $T=634260 729240 0 180 $X=633020 $Y=723820
X1070 1991 2 224 1 INV1S $T=634260 749400 1 180 $X=633020 $Y=749020
X1071 1965 2 1954 1 INV1S $T=635500 860280 1 180 $X=634260 $Y=859900
X1072 1969 2 1887 1 INV1S $T=636120 779640 1 180 $X=634880 $Y=779260
X1073 1959 2 1929 1 INV1S $T=636740 840120 1 180 $X=635500 $Y=839740
X1074 230 2 1967 1 INV1S $T=637360 729240 0 180 $X=636120 $Y=723820
X1075 1977 2 226 1 INV1S $T=637360 739320 0 180 $X=636120 $Y=733900
X1076 1968 2 1914 1 INV1S $T=636120 870360 0 0 $X=636120 $Y=869980
X1077 1973 2 1941 1 INV1S $T=639220 830040 1 180 $X=637980 $Y=829660
X1078 1984 2 1964 1 INV1S $T=639840 799800 0 180 $X=638600 $Y=794380
X1079 2003 2 1976 1 INV1S $T=641700 809880 0 180 $X=640460 $Y=804460
X1080 1988 2 1992 1 INV1S $T=640460 840120 0 0 $X=640460 $Y=839740
X1081 2032 2 1996 1 INV1S $T=644180 749400 1 180 $X=642940 $Y=749020
X1082 2011 2 1961 1 INV1S $T=644800 850200 1 180 $X=643560 $Y=849820
X1083 1997 2 2008 1 INV1S $T=644180 870360 1 0 $X=644180 $Y=864940
X1084 2002 2 1989 1 INV1S $T=646040 769560 0 180 $X=644800 $Y=764140
X1085 2022 2 233 1 INV1S $T=646660 729240 0 180 $X=645420 $Y=723820
X1086 1987 2 241 1 INV1S $T=645420 739320 0 0 $X=645420 $Y=738940
X1087 2034 2 1985 1 INV1S $T=648520 870360 0 180 $X=647280 $Y=864940
X1088 2039 2 1990 1 INV1S $T=649760 809880 1 180 $X=648520 $Y=809500
X1089 2021 2 2009 1 INV1S $T=650380 880440 1 180 $X=649140 $Y=880060
X1090 2027 2 1970 1 INV1S $T=651000 759480 1 180 $X=649760 $Y=759100
X1091 2037 2 2016 1 INV1S $T=651000 890520 1 180 $X=649760 $Y=890140
X1092 245 2 2001 1 INV1S $T=651000 900600 0 180 $X=649760 $Y=895180
X1093 2026 2 1994 1 INV1S $T=651620 779640 1 180 $X=650380 $Y=779260
X1094 1967 2 2006 1 INV1S $T=651000 729240 1 0 $X=651000 $Y=723820
X1095 2018 2 2005 1 INV1S $T=651000 799800 1 0 $X=651000 $Y=794380
X1096 2054 2 2014 1 INV1S $T=653480 799800 0 180 $X=652240 $Y=794380
X1097 199 2 2043 1 INV1S $T=652240 870360 1 0 $X=652240 $Y=864940
X1098 2061 2 2029 1 INV1S $T=654100 840120 1 180 $X=652860 $Y=839740
X1099 2052 2 2023 1 INV1S $T=656580 830040 0 180 $X=655340 $Y=824620
X1100 2028 2 2057 1 INV1S $T=656580 769560 0 0 $X=656580 $Y=769180
X1101 2053 2 1995 1 INV1S $T=657200 840120 1 0 $X=657200 $Y=834700
X1102 2073 2 248 1 INV1S $T=659060 729240 0 180 $X=657820 $Y=723820
X1103 2111 2 2040 1 INV1S $T=660300 779640 1 180 $X=659060 $Y=779260
X1104 2058 2 2035 1 INV1S $T=659060 850200 0 0 $X=659060 $Y=849820
X1105 2030 2 2064 1 INV1S $T=659060 880440 1 0 $X=659060 $Y=875020
X1106 2072 2 2004 1 INV1S $T=661540 739320 0 180 $X=660300 $Y=733900
X1107 2088 2 2076 1 INV1S $T=664020 759480 1 180 $X=662780 $Y=759100
X1108 2086 2 2080 1 INV1S $T=664020 840120 1 180 $X=662780 $Y=839740
X1109 2091 2 2079 1 INV1S $T=665260 830040 0 180 $X=664020 $Y=824620
X1110 2081 2 2048 1 INV1S $T=664640 749400 0 0 $X=664640 $Y=749020
X1111 2065 2 2094 1 INV1S $T=665260 789720 0 0 $X=665260 $Y=789340
X1112 199 2 2107 1 INV1S $T=666500 759480 0 0 $X=666500 $Y=759100
X1113 2101 2 2077 1 INV1S $T=667740 809880 1 180 $X=666500 $Y=809500
X1114 2108 2 2066 1 INV1S $T=667740 860280 0 180 $X=666500 $Y=854860
X1115 2099 2 2047 1 INV1S $T=667120 819960 1 0 $X=667120 $Y=814540
X1116 2106 2 2097 1 INV1S $T=668980 880440 1 180 $X=667740 $Y=880060
X1117 2084 2 257 1 INV1S $T=669600 719160 1 180 $X=668360 $Y=718780
X1118 2090 2 2110 1 INV1S $T=669600 749400 0 0 $X=669600 $Y=749020
X1119 260 2 259 1 INV1S $T=670840 890520 1 180 $X=669600 $Y=890140
X1120 2103 2 2115 1 INV1S $T=673940 850200 0 180 $X=672700 $Y=844780
X1121 2128 2 2125 1 INV1S $T=674560 840120 0 180 $X=673320 $Y=834700
X1122 2109 2 2139 1 INV1S $T=673940 880440 1 0 $X=673940 $Y=875020
X1123 2136 2 2089 1 INV1S $T=674560 749400 1 0 $X=674560 $Y=743980
X1124 2146 2 2141 1 INV1S $T=677040 840120 0 180 $X=675800 $Y=834700
X1125 2130 2 2124 1 INV1S $T=678280 749400 0 180 $X=677040 $Y=743980
X1126 2148 2 2119 1 INV1S $T=678280 799800 0 180 $X=677040 $Y=794380
X1127 2149 2 2126 1 INV1S $T=680140 819960 0 180 $X=678900 $Y=814540
X1128 2163 2 2155 1 INV1S $T=680760 779640 0 180 $X=679520 $Y=774220
X1129 268 2 264 1 INV1S $T=680760 900600 0 180 $X=679520 $Y=895180
X1130 2140 2 271 1 INV1S $T=680760 749400 1 0 $X=680760 $Y=743980
X1131 2142 2 2143 1 INV1S $T=681380 729240 1 0 $X=681380 $Y=723820
X1132 2162 2 2132 1 INV1S $T=682000 769560 0 0 $X=682000 $Y=769180
X1133 2167 2 2112 1 INV1S $T=683860 830040 0 180 $X=682620 $Y=824620
X1134 2182 2 2186 1 INV1S $T=685720 809880 1 0 $X=685720 $Y=804460
X1135 2191 2 2177 1 INV1S $T=686960 819960 0 180 $X=685720 $Y=814540
X1136 2192 2 2164 1 INV1S $T=686960 880440 0 180 $X=685720 $Y=875020
X1137 2116 2 2183 1 INV1S $T=685720 890520 1 0 $X=685720 $Y=885100
X1138 2189 2 2150 1 INV1S $T=687580 860280 0 180 $X=686340 $Y=854860
X1139 2195 2 2199 1 INV1S $T=688820 729240 0 0 $X=688820 $Y=728860
X1140 2203 2 2185 1 INV1S $T=690680 759480 1 180 $X=689440 $Y=759100
X1141 2213 2 2170 1 INV1S $T=690680 779640 1 180 $X=689440 $Y=779260
X1142 2211 2 2158 1 INV1S $T=691920 739320 1 180 $X=690680 $Y=738940
X1143 2206 2 2180 1 INV1S $T=691300 840120 0 0 $X=691300 $Y=839740
X1144 2212 2 2193 1 INV1S $T=693160 759480 0 0 $X=693160 $Y=759100
X1145 2215 2 2168 1 INV1S $T=694400 890520 0 180 $X=693160 $Y=885100
X1146 2232 2 2196 1 INV1S $T=695020 870360 1 180 $X=693780 $Y=869980
X1147 278 2 281 1 INV1S $T=695020 719160 0 0 $X=695020 $Y=718780
X1148 2225 2 2210 1 INV1S $T=696260 880440 0 180 $X=695020 $Y=875020
X1149 2229 2 2220 1 INV1S $T=697500 799800 1 180 $X=696260 $Y=799420
X1150 2226 2 2222 1 INV1S $T=696880 729240 0 0 $X=696880 $Y=728860
X1151 2228 2 2181 1 INV1S $T=697500 880440 1 0 $X=697500 $Y=875020
X1152 2216 2 2144 1 INV1S $T=698740 830040 0 0 $X=698740 $Y=829660
X1153 2246 2 2231 1 INV1S $T=701220 850200 1 180 $X=699980 $Y=849820
X1154 2233 2 2178 1 INV1S $T=699980 860280 0 0 $X=699980 $Y=859900
X1155 2253 2 2224 1 INV1S $T=702460 830040 1 180 $X=701220 $Y=829660
X1156 2239 2 2214 1 INV1S $T=701840 819960 1 0 $X=701840 $Y=814540
X1157 2261 2 2230 1 INV1S $T=705560 789720 1 180 $X=704320 $Y=789340
X1158 2262 2 2171 1 INV1S $T=704940 819960 1 0 $X=704940 $Y=814540
X1159 2241 2 2240 1 INV1S $T=704940 890520 1 0 $X=704940 $Y=885100
X1160 2296 2 2278 1 INV1S $T=713620 860280 1 0 $X=713620 $Y=854860
X1161 2302 2 2289 1 INV1S $T=714240 799800 0 0 $X=714240 $Y=799420
X1162 2304 2 2268 1 INV1S $T=715480 850200 1 0 $X=715480 $Y=844780
X1163 2290 2 2301 1 INV1S $T=716100 729240 0 0 $X=716100 $Y=728860
X1164 2313 2 2305 1 INV1S $T=717340 749400 0 180 $X=716100 $Y=743980
X1165 2311 2 2316 1 INV1S $T=716100 749400 0 0 $X=716100 $Y=749020
X1166 2310 2 2264 1 INV1S $T=717960 830040 0 0 $X=717960 $Y=829660
X1167 2321 2 2251 1 INV1S $T=719200 880440 1 180 $X=717960 $Y=880060
X1168 289 2 2331 1 INV1S $T=718580 739320 1 0 $X=718580 $Y=733900
X1169 2276 2 2329 1 INV1S $T=718580 749400 1 0 $X=718580 $Y=743980
X1170 2326 2 2294 1 INV1S $T=719820 850200 0 180 $X=718580 $Y=844780
X1171 2298 2 2328 1 INV1S $T=719200 759480 1 0 $X=719200 $Y=754060
X1172 2309 2 2269 1 INV1S $T=719200 830040 1 0 $X=719200 $Y=824620
X1173 2287 2 2308 1 INV1S $T=719200 870360 0 0 $X=719200 $Y=869980
X1174 2262 2 301 1 INV1S $T=719200 900600 1 0 $X=719200 $Y=895180
X1175 2325 2 2306 1 INV1S $T=719820 819960 0 0 $X=719820 $Y=819580
X1176 220 2 2262 1 INV1S $T=720440 880440 0 0 $X=720440 $Y=880060
X1177 2262 2 2236 1 INV1S $T=721060 860280 0 0 $X=721060 $Y=859900
X1178 2262 2 2344 1 INV1S $T=722300 819960 1 0 $X=722300 $Y=814540
X1179 2223 2 2334 1 INV1S $T=724780 729240 0 0 $X=724780 $Y=728860
X1180 2352 2 2345 1 INV1S $T=726640 819960 0 180 $X=725400 $Y=814540
X1181 306 2 300 1 INV1S $T=725400 900600 1 0 $X=725400 $Y=895180
X1182 2358 2 2281 1 INV1S $T=727260 890520 1 180 $X=726020 $Y=890140
X1183 2364 2 2351 1 INV1S $T=729740 870360 1 180 $X=728500 $Y=869980
X1184 2361 2 2299 1 INV1S $T=730360 809880 1 0 $X=730360 $Y=804460
X1185 2366 2 2359 1 INV1S $T=730360 850200 0 0 $X=730360 $Y=849820
X1186 2371 2 2295 1 INV1S $T=731600 890520 1 0 $X=731600 $Y=885100
X1187 2372 2 2307 1 INV1S $T=733460 870360 0 180 $X=732220 $Y=864940
X1188 2400 2 2380 1 INV1S $T=737180 739320 0 180 $X=735940 $Y=733900
X1189 322 2 2386 1 INV1S $T=739040 729240 0 180 $X=737800 $Y=723820
X1190 329 2 2385 1 INV1S $T=739660 739320 1 180 $X=738420 $Y=738940
X1191 2390 2 2350 1 INV1S $T=739040 830040 0 0 $X=739040 $Y=829660
X1192 2384 2 2409 1 INV1S $T=739040 870360 1 0 $X=739040 $Y=864940
X1193 2413 2 2363 1 INV1S $T=741520 860280 1 180 $X=740280 $Y=859900
X1194 2412 2 2379 1 INV1S $T=740900 840120 1 0 $X=740900 $Y=834700
X1195 2263 2 2408 1 INV1S $T=741520 729240 0 0 $X=741520 $Y=728860
X1196 2420 2 2399 1 INV1S $T=743380 850200 1 180 $X=742140 $Y=849820
X1197 333 2 335 1 INV1S $T=744000 719160 0 0 $X=744000 $Y=718780
X1198 2392 2 2438 1 INV1S $T=745240 890520 0 0 $X=745240 $Y=890140
X1199 2407 2 2459 1 INV1S $T=747720 769560 0 0 $X=747720 $Y=769180
X1200 2457 2 2426 1 INV1S $T=749580 799800 1 180 $X=748340 $Y=799420
X1201 2452 2 2405 1 INV1S $T=749580 830040 1 0 $X=749580 $Y=824620
X1202 2468 2 2436 1 INV1S $T=752060 830040 0 180 $X=750820 $Y=824620
X1203 325 2 2474 1 INV1S $T=751440 799800 0 0 $X=751440 $Y=799420
X1204 2476 2 2444 1 INV1S $T=753300 850200 0 180 $X=752060 $Y=844780
X1205 2454 2 2482 1 INV1S $T=753300 779640 0 0 $X=753300 $Y=779260
X1206 2466 2 2463 1 INV1S $T=753920 850200 0 0 $X=753920 $Y=849820
X1207 2472 2 339 1 INV1S $T=753920 870360 1 0 $X=753920 $Y=864940
X1208 2467 2 2490 1 INV1S $T=755160 749400 0 0 $X=755160 $Y=749020
X1209 2447 2 2495 1 INV1S $T=755780 779640 0 0 $X=755780 $Y=779260
X1210 2330 2 346 1 INV1S $T=756400 719160 0 0 $X=756400 $Y=718780
X1211 343 2 2496 1 INV1S $T=756400 729240 1 0 $X=756400 $Y=723820
X1212 2503 2 2465 1 INV1S $T=758260 739320 0 180 $X=757020 $Y=733900
X1213 2488 2 2464 1 INV1S $T=757020 860280 1 0 $X=757020 $Y=854860
X1214 344 2 2503 1 INV1S $T=758880 729240 1 180 $X=757640 $Y=728860
X1215 2510 2 2497 1 INV1S $T=759500 830040 0 180 $X=758260 $Y=824620
X1216 2503 2 2516 1 INV1S $T=758880 739320 1 0 $X=758880 $Y=733900
X1217 2471 2 2505 1 INV1S $T=760120 759480 1 0 $X=760120 $Y=754060
X1218 2517 2 2483 1 INV1S $T=760120 809880 0 0 $X=760120 $Y=809500
X1219 2439 2 2521 1 INV1S $T=760740 739320 0 0 $X=760740 $Y=738940
X1220 349 2 2512 1 INV1S $T=761980 900600 0 180 $X=760740 $Y=895180
X1221 2416 2 2509 1 INV1S $T=761360 759480 1 0 $X=761360 $Y=754060
X1222 2518 2 2492 1 INV1S $T=761980 890520 0 0 $X=761980 $Y=890140
X1223 2529 2 2535 1 INV1S $T=762600 749400 0 0 $X=762600 $Y=749020
X1224 2501 2 2525 1 INV1S $T=762600 880440 0 0 $X=762600 $Y=880060
X1225 2489 2 2528 1 INV1S $T=763840 729240 1 0 $X=763840 $Y=723820
X1226 2543 2 2504 1 INV1S $T=765080 799800 0 180 $X=763840 $Y=794380
X1227 2565 2 2491 1 INV1S $T=765080 840120 1 180 $X=763840 $Y=839740
X1228 2546 2 2500 1 INV1S $T=765080 860280 1 180 $X=763840 $Y=859900
X1229 2489 2 2549 1 INV1S $T=764460 719160 0 0 $X=764460 $Y=718780
X1230 2456 2 2557 1 INV1S $T=766320 789720 1 0 $X=766320 $Y=784300
X1231 2542 2 2544 1 INV1S $T=766940 799800 0 0 $X=766940 $Y=799420
X1232 2558 2 2546 1 INV1S $T=766940 870360 0 0 $X=766940 $Y=869980
X1233 2560 2 2573 1 INV1S $T=768800 769560 1 0 $X=768800 $Y=764140
X1234 2383 2 2569 1 INV1S $T=768800 809880 0 0 $X=768800 $Y=809500
X1235 210 2 2558 1 INV1S $T=768800 900600 1 0 $X=768800 $Y=895180
X1236 2577 2 2530 1 INV1S $T=771280 819960 1 180 $X=770040 $Y=819580
X1237 2540 2 2584 1 INV1S $T=770660 769560 0 0 $X=770660 $Y=769180
X1238 2582 2 2548 1 INV1S $T=771900 809880 1 180 $X=770660 $Y=809500
X1239 2283 2 2581 1 INV1S $T=771900 739320 1 0 $X=771900 $Y=733900
X1240 2297 2 2605 1 INV1S $T=775620 729240 1 0 $X=775620 $Y=723820
X1241 2596 2 356 1 INV1S $T=775620 880440 0 0 $X=775620 $Y=880060
X1242 2502 2 2594 1 INV1S $T=776240 779640 0 0 $X=776240 $Y=779260
X1243 2606 2 2595 1 INV1S $T=777480 799800 1 180 $X=776240 $Y=799420
X1244 2608 2 358 1 INV1S $T=777480 890520 1 180 $X=776240 $Y=890140
X1245 2576 2 2629 1 INV1S $T=779340 799800 1 0 $X=779340 $Y=794380
X1246 113 2 2619 1 INV1S $T=781200 819960 0 180 $X=779960 $Y=814540
X1247 2617 2 2593 1 INV1S $T=781200 860280 0 0 $X=781200 $Y=859900
X1248 2614 2 2627 1 INV1S $T=784920 779640 0 180 $X=783680 $Y=774220
X1249 2637 2 2570 1 INV1S $T=784920 860280 1 180 $X=783680 $Y=859900
X1250 2633 2 2640 1 INV1S $T=784300 759480 1 0 $X=784300 $Y=754060
X1251 2644 2 2591 1 INV1S $T=786780 850200 1 180 $X=785540 $Y=849820
X1252 2654 2 2634 1 INV1S $T=788020 840120 1 180 $X=786780 $Y=839740
X1253 2645 2 367 1 INV1S $T=786780 870360 0 0 $X=786780 $Y=869980
X1254 2657 2 2626 1 INV1S $T=788640 830040 0 180 $X=787400 $Y=824620
X1255 2639 2 2662 1 INV1S $T=789260 759480 1 0 $X=789260 $Y=754060
X1256 2668 2 362 1 INV1S $T=791120 880440 1 180 $X=789880 $Y=880060
X1257 2673 2 2620 1 INV1S $T=792360 809880 1 180 $X=791120 $Y=809500
X1258 2288 2 2675 1 INV1S $T=791740 729240 1 0 $X=791740 $Y=723820
X1259 2698 2 370 1 INV1S $T=794220 870360 0 180 $X=792980 $Y=864940
X1260 2684 2 2672 1 INV1S $T=794840 799800 1 180 $X=793600 $Y=799420
X1261 364 2 2706 1 INV1S $T=794220 900600 1 0 $X=794220 $Y=895180
X1262 2688 2 372 1 INV1S $T=796080 850200 1 180 $X=794840 $Y=849820
X1263 2674 2 2693 1 INV1S $T=795460 739320 1 0 $X=795460 $Y=733900
X1264 2651 2 2690 1 INV1S $T=795460 759480 0 0 $X=795460 $Y=759100
X1265 2664 2 2700 1 INV1S $T=796080 739320 0 0 $X=796080 $Y=738940
X1266 2647 2 2692 1 INV1S $T=796080 759480 1 0 $X=796080 $Y=754060
X1267 2699 2 374 1 INV1S $T=797940 870360 0 0 $X=797940 $Y=869980
X1268 2721 2 371 1 INV1S $T=799180 890520 1 180 $X=797940 $Y=890140
X1269 2703 2 382 1 INV1S $T=800420 860280 0 0 $X=800420 $Y=859900
X1270 2725 2 2686 1 INV1S $T=804140 830040 0 180 $X=802900 $Y=824620
X1271 2734 2 2717 1 INV1S $T=806000 830040 1 180 $X=804760 $Y=829660
X1272 386 2 379 1 INV1S $T=806620 890520 1 180 $X=805380 $Y=890140
X1273 2753 2 2708 1 INV1S $T=807860 819960 0 180 $X=806620 $Y=814540
X1274 2737 2 2694 1 INV1S $T=808480 840120 0 180 $X=807240 $Y=834700
X1275 2754 2 384 1 INV1S $T=809100 840120 1 180 $X=807860 $Y=839740
X1276 2757 2 377 1 INV1S $T=812820 860280 0 180 $X=811580 $Y=854860
X1277 2706 2 393 1 INV1S $T=814060 900600 1 0 $X=814060 $Y=895180
X1278 2759 2 387 1 INV1S $T=815920 870360 0 180 $X=814680 $Y=864940
X1279 2752 2 390 1 INV1S $T=814680 880440 0 0 $X=814680 $Y=880060
X1280 2658 2 2761 1 INV1S $T=815920 739320 0 0 $X=815920 $Y=738940
X1281 2778 2 389 1 INV1S $T=817160 870360 0 180 $X=815920 $Y=864940
X1282 2785 2 388 1 INV1S $T=819020 880440 1 180 $X=817780 $Y=880060
X1283 2779 2 2775 1 INV1S $T=820880 729240 0 180 $X=819640 $Y=723820
X1284 2787 2 2764 1 INV1S $T=821500 840120 1 180 $X=820260 $Y=839740
X1285 2784 2 2782 1 INV1S $T=822740 719160 1 180 $X=821500 $Y=718780
X1286 2788 2 2795 1 INV1S $T=821500 749400 0 0 $X=821500 $Y=749020
X1287 2834 2 2818 1 INV1S $T=828940 749400 1 180 $X=827700 $Y=749020
X1288 2814 2 2835 1 INV1S $T=828320 870360 0 0 $X=828320 $Y=869980
X1289 2815 2 403 1 INV1S $T=829560 719160 0 0 $X=829560 $Y=718780
X1290 2846 2 2830 1 INV1S $T=830800 860280 1 180 $X=829560 $Y=859900
X1291 2824 2 2839 1 INV1S $T=831420 870360 1 180 $X=830180 $Y=869980
X1292 2850 2 2829 1 INV1S $T=832040 799800 0 180 $X=830800 $Y=794380
X1293 2864 2 2842 1 INV1S $T=832040 860280 1 180 $X=830800 $Y=859900
X1294 2801 2 2836 1 INV1S $T=832040 890520 0 180 $X=830800 $Y=885100
X1295 2860 2 2828 1 INV1S $T=832660 779640 1 180 $X=831420 $Y=779260
X1296 2853 2 2866 1 INV1S $T=832660 860280 1 0 $X=832660 $Y=854860
X1297 2869 2 2858 1 INV1S $T=833900 870360 1 180 $X=832660 $Y=869980
X1298 2841 2 2859 1 INV1S $T=834520 819960 1 180 $X=833280 $Y=819580
X1299 2855 2 2871 1 INV1S $T=833900 749400 1 0 $X=833900 $Y=743980
X1300 2867 2 2845 1 INV1S $T=834520 779640 1 0 $X=834520 $Y=774220
X1301 2872 2 2881 1 INV1S $T=836380 739320 0 0 $X=836380 $Y=738940
X1302 2857 2 2865 1 INV1S $T=838240 809880 0 180 $X=837000 $Y=804460
X1303 2800 2 2886 1 INV1S $T=840100 830040 1 0 $X=840100 $Y=824620
X1304 2892 2 2904 1 INV1S $T=841960 850200 0 0 $X=841960 $Y=849820
X1305 2895 2 2907 1 INV1S $T=843200 870360 1 0 $X=843200 $Y=864940
X1306 2910 2 2908 1 INV1S $T=846920 819960 0 180 $X=845680 $Y=814540
X1307 2921 2 2894 1 INV1S $T=847540 789720 1 180 $X=846300 $Y=789340
X1308 398 2 2900 1 INV1S $T=848780 890520 1 180 $X=847540 $Y=890140
X1309 2940 2 2933 1 INV1S $T=850640 850200 1 180 $X=849400 $Y=849820
X1310 2918 2 2951 1 INV1S $T=850020 880440 1 0 $X=850020 $Y=875020
X1311 2948 2 2956 1 INV1S $T=850640 749400 1 0 $X=850640 $Y=743980
X1312 2912 2 2955 1 INV1S $T=851260 819960 0 0 $X=851260 $Y=819580
X1313 2957 2 2943 1 INV1S $T=853120 769560 1 180 $X=851880 $Y=769180
X1314 2939 2 2883 1 INV1S $T=853120 799800 0 180 $X=851880 $Y=794380
X1315 2936 2 2942 1 INV1S $T=853740 759480 0 180 $X=852500 $Y=754060
X1316 2968 2 2944 1 INV1S $T=853740 779640 0 180 $X=852500 $Y=774220
X1317 2964 2 2959 1 INV1S $T=854360 759480 1 180 $X=853120 $Y=759100
X1318 2975 2 2954 1 INV1S $T=855600 809880 0 180 $X=854360 $Y=804460
X1319 428 2 2990 1 INV1S $T=855600 870360 1 0 $X=855600 $Y=864940
X1320 2988 2 2963 1 INV1S $T=857460 870360 1 180 $X=856220 $Y=869980
X1321 2986 2 2960 1 INV1S $T=858080 749400 1 180 $X=856840 $Y=749020
X1322 2995 2 2977 1 INV1S $T=859320 739320 1 180 $X=858080 $Y=738940
X1323 2949 2 2966 1 INV1S $T=859320 890520 0 180 $X=858080 $Y=885100
X1324 2980 2 2931 1 INV1S $T=859940 779640 0 180 $X=858700 $Y=774220
X1325 2973 2 3004 1 INV1S $T=858700 809880 1 0 $X=858700 $Y=804460
X1326 2985 2 2983 1 INV1S $T=859940 850200 1 180 $X=858700 $Y=849820
X1327 2938 2 2979 1 INV1S $T=860560 860280 1 180 $X=859320 $Y=859900
X1328 2992 2 2998 1 INV1S $T=861800 769560 0 180 $X=860560 $Y=764140
X1329 2923 2 2993 1 INV1S $T=861800 840120 0 0 $X=861800 $Y=839740
X1330 3008 2 3030 1 INV1S $T=863040 769560 1 0 $X=863040 $Y=764140
X1331 3042 2 2938 1 INV1S $T=864900 870360 0 180 $X=863660 $Y=864940
X1332 3007 2 2999 1 INV1S $T=866140 830040 1 180 $X=864900 $Y=829660
X1333 3021 2 3045 1 INV1S $T=865520 779640 1 0 $X=865520 $Y=774220
X1334 3042 2 2976 1 INV1S $T=868000 870360 0 180 $X=866760 $Y=864940
X1335 3053 2 3011 1 INV1S $T=869240 729240 0 180 $X=868000 $Y=723820
X1336 3102 2 3024 1 INV1S $T=869860 809880 0 180 $X=868620 $Y=804460
X1337 3068 2 3036 1 INV1S $T=870480 749400 1 180 $X=869240 $Y=749020
X1338 3060 2 3050 1 INV1S $T=871100 870360 1 180 $X=869860 $Y=869980
X1339 3018 2 3052 1 INV1S $T=871720 759480 1 180 $X=870480 $Y=759100
X1340 3065 2 3088 1 INV1S $T=871720 860280 0 0 $X=871720 $Y=859900
X1341 448 2 443 1 INV1S $T=873580 890520 1 180 $X=872340 $Y=890140
X1342 3087 2 3061 1 INV1S $T=874200 779640 0 180 $X=872960 $Y=774220
X1343 3009 2 426 1 INV1S $T=874200 870360 1 180 $X=872960 $Y=869980
X1344 3099 2 3085 1 INV1S $T=875440 749400 1 180 $X=874200 $Y=749020
X1345 3080 2 3096 1 INV1S $T=877300 809880 1 180 $X=876060 $Y=809500
X1346 3042 2 3079 1 INV1S $T=876060 870360 1 0 $X=876060 $Y=864940
X1347 3086 2 3095 1 INV1S $T=877920 769560 0 180 $X=876680 $Y=764140
X1348 3067 2 3116 1 INV1S $T=877300 900600 1 0 $X=877300 $Y=895180
X1349 3103 2 3122 1 INV1S $T=878540 789720 1 0 $X=878540 $Y=784300
X1350 3070 2 3128 1 INV1S $T=879160 819960 1 0 $X=879160 $Y=814540
X1351 3075 2 3083 1 INV1S $T=879780 749400 0 0 $X=879780 $Y=749020
X1352 3142 2 3043 1 INV1S $T=883500 799800 1 0 $X=883500 $Y=794380
X1353 3121 2 3132 1 INV1S $T=885360 749400 1 0 $X=885360 $Y=743980
X1354 3167 2 3164 1 INV1S $T=887840 880440 0 180 $X=886600 $Y=875020
X1355 3169 2 3150 1 INV1S $T=889080 749400 0 180 $X=887840 $Y=743980
X1356 3153 2 3188 1 INV1S $T=889700 769560 1 0 $X=889700 $Y=764140
X1357 3133 2 3182 1 INV1S $T=891560 769560 1 180 $X=890320 $Y=769180
X1358 3201 2 3135 1 INV1S $T=894040 809880 1 180 $X=892800 $Y=809500
X1359 3185 2 3213 1 INV1S $T=892800 840120 0 0 $X=892800 $Y=839740
X1360 3148 2 3211 1 INV1S $T=892800 860280 0 0 $X=892800 $Y=859900
X1361 3184 2 3192 1 INV1S $T=893420 860280 1 0 $X=893420 $Y=854860
X1362 3205 2 3217 1 INV1S $T=894660 830040 1 0 $X=894660 $Y=824620
X1363 3199 2 3189 1 INV1S $T=895280 830040 0 0 $X=895280 $Y=829660
X1364 3209 2 3222 1 INV1S $T=895280 880440 1 0 $X=895280 $Y=875020
X1365 3196 2 3232 1 INV1S $T=895900 789720 0 0 $X=895900 $Y=789340
X1366 3214 2 3238 1 INV1S $T=896520 729240 0 0 $X=896520 $Y=728860
X1367 3198 2 3172 1 INV1S $T=896520 759480 0 0 $X=896520 $Y=759100
X1368 3151 2 3223 1 INV1S $T=896520 850200 1 0 $X=896520 $Y=844780
X1369 3086 2 3229 1 INV1S $T=897140 749400 0 0 $X=897140 $Y=749020
X1370 3212 2 3227 1 INV1S $T=899000 719160 0 0 $X=899000 $Y=718780
X1371 3069 2 3005 1 INV1S $T=899620 749400 1 0 $X=899620 $Y=743980
X1372 3220 2 3259 1 INV1S $T=900860 739320 1 0 $X=900860 $Y=733900
X1373 3260 2 3156 1 INV1S $T=902720 759480 1 180 $X=901480 $Y=759100
X1374 482 2 3262 1 INV1S $T=902100 870360 1 0 $X=902100 $Y=864940
X1375 2683 2 3249 1 INV1S $T=902720 779640 0 0 $X=902720 $Y=779260
X1376 3275 2 3266 1 INV1S $T=904580 880440 0 180 $X=903340 $Y=875020
X1377 2792 2 3163 1 INV1S $T=903960 789720 1 0 $X=903960 $Y=784300
X1378 3251 2 3269 1 INV1S $T=903960 830040 0 0 $X=903960 $Y=829660
X1379 3174 2 3260 1 INV1S $T=905200 769560 1 0 $X=905200 $Y=764140
X1380 3288 2 3248 1 INV1S $T=907060 759480 1 180 $X=905820 $Y=759100
X1381 3264 2 3291 1 INV1S $T=905820 880440 0 0 $X=905820 $Y=880060
X1382 3193 2 3290 1 INV1S $T=906440 850200 1 0 $X=906440 $Y=844780
X1383 3243 2 3300 1 INV1S $T=907680 850200 0 0 $X=907680 $Y=849820
X1384 461 2 486 1 INV1S $T=907680 900600 1 0 $X=907680 $Y=895180
X1385 3256 2 3286 1 INV1S $T=908300 729240 1 0 $X=908300 $Y=723820
X1386 3260 2 3316 1 INV1S $T=908300 769560 1 0 $X=908300 $Y=764140
X1387 3287 2 3312 1 INV1S $T=908920 729240 0 0 $X=908920 $Y=728860
X1388 3289 2 3309 1 INV1S $T=910160 779640 0 0 $X=910160 $Y=779260
X1389 3295 2 487 1 INV1S $T=910780 719160 0 0 $X=910780 $Y=718780
X1390 3225 2 3315 1 INV1S $T=910780 880440 1 0 $X=910780 $Y=875020
X1391 3304 2 489 1 INV1S $T=912020 719160 0 0 $X=912020 $Y=718780
X1392 3323 2 3326 1 INV1S $T=912020 759480 1 0 $X=912020 $Y=754060
X1393 3317 2 3268 1 INV1S $T=912020 779640 1 0 $X=912020 $Y=774220
X1394 3329 2 3349 1 INV1S $T=916360 739320 0 0 $X=916360 $Y=738940
X1395 3311 2 3336 1 INV1S $T=916360 830040 0 0 $X=916360 $Y=829660
X1396 3347 2 3376 1 INV1S $T=918840 830040 0 0 $X=918840 $Y=829660
X1397 3360 2 3362 1 INV1S $T=920700 729240 0 180 $X=919460 $Y=723820
X1398 3383 2 3301 1 INV1S $T=922560 799800 1 180 $X=921320 $Y=799420
X1399 3384 2 3382 1 INV1S $T=923800 759480 0 180 $X=922560 $Y=754060
X1400 3334 2 3389 1 INV1S $T=923180 860280 1 0 $X=923180 $Y=854860
X1401 3278 2 3391 1 INV1S $T=923180 900600 1 0 $X=923180 $Y=895180
X1402 3365 2 3403 1 INV1S $T=924420 860280 1 0 $X=924420 $Y=854860
X1403 3276 2 3346 1 INV1S $T=925040 779640 0 0 $X=925040 $Y=779260
X1404 3371 2 3394 1 INV1S $T=925040 850200 1 0 $X=925040 $Y=844780
X1405 2741 2 3407 1 INV1S $T=926900 789720 1 0 $X=926900 $Y=784300
X1406 3399 2 3386 1 INV1S $T=927520 719160 0 0 $X=927520 $Y=718780
X1407 3412 2 3419 1 INV1S $T=928760 739320 0 0 $X=928760 $Y=738940
X1408 3388 2 3438 1 INV1S $T=929380 799800 1 0 $X=929380 $Y=794380
X1409 3405 2 3422 1 INV1S $T=930000 759480 1 0 $X=930000 $Y=754060
X1410 3423 2 3374 1 INV1S $T=931240 769560 1 180 $X=930000 $Y=769180
X1411 3366 2 3435 1 INV1S $T=931240 789720 0 0 $X=931240 $Y=789340
X1412 3388 2 3409 1 INV1S $T=933720 789720 0 180 $X=932480 $Y=784300
X1413 3426 2 3439 1 INV1S $T=932480 850200 0 0 $X=932480 $Y=849820
X1414 3398 2 3441 1 INV1S $T=932480 870360 0 0 $X=932480 $Y=869980
X1415 3121 2 3452 1 INV1S $T=933720 749400 0 0 $X=933720 $Y=749020
X1416 3397 2 3450 1 INV1S $T=934340 729240 0 0 $X=934340 $Y=728860
X1417 3121 2 3468 1 INV1S $T=934960 739320 1 0 $X=934960 $Y=733900
X1418 3388 2 3456 1 INV1S $T=934960 789720 1 0 $X=934960 $Y=784300
X1419 3388 2 3445 1 INV1S $T=934960 799800 0 0 $X=934960 $Y=799420
X1420 3406 2 3454 1 INV1S $T=935580 850200 0 0 $X=935580 $Y=849820
X1421 3447 2 3473 1 INV1S $T=938060 759480 1 0 $X=938060 $Y=754060
X1422 3465 2 3485 1 INV1S $T=939300 729240 1 0 $X=939300 $Y=723820
X1423 3265 2 3451 1 INV1S $T=939300 749400 0 0 $X=939300 $Y=749020
X1424 3408 2 3471 1 INV1S $T=941780 779640 0 180 $X=940540 $Y=774220
X1425 3434 2 3482 1 INV1S $T=940540 880440 1 0 $X=940540 $Y=875020
X1426 3481 2 3497 1 INV1S $T=942400 850200 1 0 $X=942400 $Y=844780
X1427 3476 2 3495 1 INV1S $T=943020 789720 1 0 $X=943020 $Y=784300
X1428 3480 2 3489 1 INV1S $T=944880 759480 1 180 $X=943640 $Y=759100
X1429 3499 2 3494 1 INV1S $T=944880 860280 1 180 $X=943640 $Y=859900
X1430 521 2 3500 1 INV1S $T=944260 729240 0 0 $X=944260 $Y=728860
X1431 3421 2 3505 1 INV1S $T=944260 739320 0 0 $X=944260 $Y=738940
X1432 3402 2 3511 1 INV1S $T=944880 789720 0 0 $X=944880 $Y=789340
X1433 3483 2 3509 1 INV1S $T=951080 850200 1 0 $X=951080 $Y=844780
X1434 3525 2 3539 1 INV1S $T=951700 799800 1 0 $X=951700 $Y=794380
X1435 535 2 3540 1 INV1S $T=951700 890520 1 0 $X=951700 $Y=885100
X1436 3487 2 3541 1 INV1S $T=953560 840120 0 0 $X=953560 $Y=839740
X1437 537 2 3550 1 INV1S $T=955420 890520 1 180 $X=954180 $Y=890140
X1438 3516 2 3549 1 INV1S $T=956040 779640 0 0 $X=956040 $Y=779260
X1439 3546 2 3529 1 INV1S $T=956040 880440 0 0 $X=956040 $Y=880060
X1440 3501 2 3559 1 INV1S $T=957280 769560 1 0 $X=957280 $Y=764140
X1441 3520 2 3552 1 INV1S $T=958520 799800 1 0 $X=958520 $Y=794380
X1442 3532 2 3571 1 INV1S $T=959760 759480 0 0 $X=959760 $Y=759100
X1443 3563 2 3572 1 INV1S $T=960380 739320 0 0 $X=960380 $Y=738940
X1444 3570 2 3588 1 INV1S $T=962240 749400 1 0 $X=962240 $Y=743980
X1445 3536 2 3586 1 INV1S $T=962860 759480 1 0 $X=962860 $Y=754060
X1446 3565 2 3598 1 INV1S $T=963480 739320 1 0 $X=963480 $Y=733900
X1447 3562 2 3602 1 INV1S $T=967200 769560 1 0 $X=967200 $Y=764140
X1448 3555 2 3607 1 INV1S $T=967820 739320 1 0 $X=967820 $Y=733900
X1449 3436 2 3584 1 INV1S $T=970920 799800 0 0 $X=970920 $Y=799420
X1450 550 2 3629 1 INV1S $T=971540 900600 1 0 $X=971540 $Y=895180
X1451 3493 2 3633 1 INV1S $T=976500 779640 1 0 $X=976500 $Y=774220
X1452 556 2 3641 1 INV1S $T=985180 719160 1 180 $X=983940 $Y=718780
X1453 3616 2 3648 1 INV1S $T=987040 779640 1 0 $X=987040 $Y=774220
X1454 3650 2 3636 1 INV1S $T=989520 749400 0 0 $X=989520 $Y=749020
X1455 611 606 591 598 2 1 MXL2HS $T=317440 789720 0 180 $X=311860 $Y=784300
X1456 660 655 630 643 2 1 MXL2HS $T=332320 779640 1 180 $X=326740 $Y=779260
X1457 29 28 25 771 2 1 MXL2HS $T=367660 900600 0 180 $X=362080 $Y=895180
X1458 771 28 802 807 2 1 MXL2HS $T=365800 890520 0 0 $X=365800 $Y=890140
X1459 807 28 792 836 2 1 MXL2HS $T=373240 880440 0 0 $X=373240 $Y=880060
X1460 35 28 33 823 2 1 MXL2HS $T=379440 900600 0 180 $X=373860 $Y=895180
X1461 823 28 809 848 2 1 MXL2HS $T=375100 890520 0 0 $X=375100 $Y=890140
X1462 847 858 814 876 2 1 MXL2HS $T=380060 870360 0 0 $X=380060 $Y=869980
X1463 836 858 796 877 2 1 MXL2HS $T=380060 880440 1 0 $X=380060 $Y=875020
X1464 880 858 865 847 2 1 MXL2HS $T=386260 880440 1 180 $X=380680 $Y=880060
X1465 885 883 839 867 2 1 MXL2HS $T=387500 850200 0 180 $X=381920 $Y=844780
X1466 848 42 890 900 2 1 MXL2HS $T=383780 890520 1 0 $X=383780 $Y=885100
X1467 43 42 896 880 2 1 MXL2HS $T=384400 890520 0 0 $X=384400 $Y=890140
X1468 877 883 808 885 2 1 MXL2HS $T=391840 860280 1 180 $X=386260 $Y=859900
X1469 867 914 922 931 2 1 MXL2HS $T=391840 840120 1 0 $X=391840 $Y=834700
X1470 876 883 927 932 2 1 MXL2HS $T=391840 860280 0 0 $X=391840 $Y=859900
X1471 932 883 895 916 2 1 MXL2HS $T=398040 850200 0 180 $X=392460 $Y=844780
X1472 900 858 957 966 2 1 MXL2HS $T=399280 880440 1 0 $X=399280 $Y=875020
X1473 951 914 947 969 2 1 MXL2HS $T=399900 840120 1 0 $X=399900 $Y=834700
X1474 916 914 874 951 2 1 MXL2HS $T=400520 840120 0 0 $X=400520 $Y=839740
X1475 966 971 964 990 2 1 MXL2HS $T=403620 870360 1 0 $X=403620 $Y=864940
X1476 931 984 919 1005 2 1 MXL2HS $T=406100 830040 1 0 $X=406100 $Y=824620
X1477 969 984 997 1010 2 1 MXL2HS $T=406720 819960 0 0 $X=406720 $Y=819580
X1478 990 971 956 1014 2 1 MXL2HS $T=407340 860280 0 0 $X=407340 $Y=859900
X1479 1005 984 1016 1037 2 1 MXL2HS $T=414160 819960 0 0 $X=414160 $Y=819580
X1480 1042 64 995 1030 2 1 MXL2HS $T=420980 880440 1 180 $X=415400 $Y=880060
X1481 1053 971 1027 1038 2 1 MXL2HS $T=423460 860280 1 180 $X=417880 $Y=859900
X1482 1030 64 1028 1053 2 1 MXL2HS $T=417880 880440 1 0 $X=417880 $Y=875020
X1483 65 64 972 1042 2 1 MXL2HS $T=424700 900600 0 180 $X=419120 $Y=895180
X1484 1047 1048 1058 1063 2 1 MXL2HS $T=419740 830040 0 0 $X=419740 $Y=829660
X1485 1038 971 1055 1047 2 1 MXL2HS $T=419740 850200 0 0 $X=419740 $Y=849820
X1486 1014 971 948 1080 2 1 MXL2HS $T=425320 850200 0 0 $X=425320 $Y=849820
X1487 1063 1048 1064 1077 2 1 MXL2HS $T=426560 830040 0 0 $X=426560 $Y=829660
X1488 1010 1074 1057 1087 2 1 MXL2HS $T=427180 819960 1 0 $X=427180 $Y=814540
X1489 1077 1048 1060 1089 2 1 MXL2HS $T=428420 819960 0 0 $X=428420 $Y=819580
X1490 74 76 1061 1091 2 1 MXL2HS $T=428420 890520 1 0 $X=428420 $Y=885100
X1491 1037 1074 1096 1113 2 1 MXL2HS $T=432760 819960 1 0 $X=432760 $Y=814540
X1492 1087 1110 1095 1124 2 1 MXL2HS $T=435240 799800 0 0 $X=435240 $Y=799420
X1493 1112 1048 1120 1128 2 1 MXL2HS $T=435860 830040 0 0 $X=435860 $Y=829660
X1494 1116 1129 1085 1115 2 1 MXL2HS $T=442680 870360 1 180 $X=437100 $Y=869980
X1495 1091 1130 1107 1116 2 1 MXL2HS $T=442680 880440 1 180 $X=437100 $Y=880060
X1496 1080 1126 1111 1112 2 1 MXL2HS $T=438960 850200 1 0 $X=438960 $Y=844780
X1497 1128 1110 1135 1134 2 1 MXL2HS $T=440200 819960 0 0 $X=440200 $Y=819580
X1498 1123 1129 1138 1143 2 1 MXL2HS $T=440200 860280 0 0 $X=440200 $Y=859900
X1499 1134 1110 1118 1145 2 1 MXL2HS $T=441440 799800 0 0 $X=441440 $Y=799420
X1500 1089 1110 1137 1149 2 1 MXL2HS $T=442680 809880 0 0 $X=442680 $Y=809500
X1501 1115 1129 1084 1123 2 1 MXL2HS $T=449500 870360 0 180 $X=443920 $Y=864940
X1502 1151 1129 1160 1162 2 1 MXL2HS $T=447020 860280 0 0 $X=447020 $Y=859900
X1503 1152 1129 1144 1151 2 1 MXL2HS $T=447020 870360 0 0 $X=447020 $Y=869980
X1504 1143 1126 1166 1174 2 1 MXL2HS $T=448880 850200 1 0 $X=448880 $Y=844780
X1505 1149 1172 1189 1184 2 1 MXL2HS $T=453840 799800 1 0 $X=453840 $Y=794380
X1506 1162 1126 1193 1195 2 1 MXL2HS $T=454460 850200 0 0 $X=454460 $Y=849820
X1507 1174 1197 1192 1185 2 1 MXL2HS $T=461280 830040 0 180 $X=455700 $Y=824620
X1508 1195 1126 1141 1203 2 1 MXL2HS $T=456940 830040 0 0 $X=456940 $Y=829660
X1509 1124 1172 1201 108 2 1 MXL2HS $T=457560 779640 0 0 $X=457560 $Y=779260
X1510 1185 1197 1196 1210 2 1 MXL2HS $T=458800 819960 1 0 $X=458800 $Y=814540
X1511 1113 1172 1208 1211 2 1 MXL2HS $T=459420 799800 1 0 $X=459420 $Y=794380
X1512 1203 1197 1217 1216 2 1 MXL2HS $T=463760 830040 1 0 $X=463760 $Y=824620
X1513 110 97 1218 1228 2 1 MXL2HS $T=463760 890520 0 0 $X=463760 $Y=890140
X1514 1145 1172 1219 112 2 1 MXL2HS $T=464380 779640 0 0 $X=464380 $Y=779260
X1515 1216 1197 1198 1236 2 1 MXL2HS $T=465620 819960 0 0 $X=465620 $Y=819580
X1516 1210 1172 1230 1235 2 1 MXL2HS $T=466240 799800 1 0 $X=466240 $Y=794380
X1517 1215 1226 1233 1240 2 1 MXL2HS $T=466860 870360 1 0 $X=466860 $Y=864940
X1518 1246 1238 1214 1229 2 1 MXL2HS $T=473680 840120 1 180 $X=468100 $Y=839740
X1519 1184 1241 1225 117 2 1 MXL2HS $T=469960 779640 1 0 $X=469960 $Y=774220
X1520 1229 1238 1232 1254 2 1 MXL2HS $T=469960 830040 1 0 $X=469960 $Y=824620
X1521 1240 1226 1221 1246 2 1 MXL2HS $T=469960 860280 0 0 $X=469960 $Y=859900
X1522 1258 1251 1212 115 2 1 MXL2HS $T=476160 759480 0 180 $X=470580 $Y=754060
X1523 1235 1241 1187 119 2 1 MXL2HS $T=470580 769560 1 0 $X=470580 $Y=764140
X1524 1211 1241 1188 120 2 1 MXL2HS $T=473060 769560 0 0 $X=473060 $Y=769180
X1525 1260 1262 1237 116 2 1 MXL2HS $T=478640 789720 0 180 $X=473060 $Y=784300
X1526 1272 1226 1239 1215 2 1 MXL2HS $T=479260 870360 0 180 $X=473680 $Y=864940
X1527 1276 121 1243 118 2 1 MXL2HS $T=479880 719160 1 180 $X=474300 $Y=718780
X1528 1228 1130 1266 1272 2 1 MXL2HS $T=474300 880440 0 0 $X=474300 $Y=880060
X1529 1254 1275 1245 1259 2 1 MXL2HS $T=480500 819960 0 180 $X=474920 $Y=814540
X1530 1280 1275 1263 1260 2 1 MXL2HS $T=480500 819960 1 180 $X=474920 $Y=819580
X1531 1285 1226 1284 1274 2 1 MXL2HS $T=483600 860280 1 180 $X=478020 $Y=859900
X1532 1305 1262 1252 1258 2 1 MXL2HS $T=484840 789720 0 180 $X=479260 $Y=784300
X1533 1307 1299 1257 1285 2 1 MXL2HS $T=484840 890520 1 180 $X=479260 $Y=890140
X1534 1271 1238 1298 1309 2 1 MXL2HS $T=479880 830040 0 0 $X=479880 $Y=829660
X1535 1297 121 1277 123 2 1 MXL2HS $T=486080 719160 1 180 $X=480500 $Y=718780
X1536 1288 1241 1269 124 2 1 MXL2HS $T=480500 769560 0 0 $X=480500 $Y=769180
X1537 1274 1238 1303 1280 2 1 MXL2HS $T=480500 840120 0 0 $X=480500 $Y=839740
X1538 1313 1251 1292 1276 2 1 MXL2HS $T=486700 759480 0 180 $X=481120 $Y=754060
X1539 1259 1293 1290 1314 2 1 MXL2HS $T=481120 799800 0 0 $X=481120 $Y=799420
X1540 1300 1282 1312 1318 2 1 MXL2HS $T=482360 779640 0 0 $X=482360 $Y=779260
X1541 1270 1251 1319 125 2 1 MXL2HS $T=482980 749400 0 0 $X=482980 $Y=749020
X1542 1316 1226 1304 1271 2 1 MXL2HS $T=489800 860280 1 180 $X=484220 $Y=859900
X1543 1329 1293 1321 1270 2 1 MXL2HS $T=491040 789720 1 180 $X=485460 $Y=789340
X1544 1318 121 1317 131 2 1 MXL2HS $T=487320 719160 0 0 $X=487320 $Y=718780
X1545 1278 1346 1332 128 2 1 MXL2HS $T=495380 729240 1 180 $X=489800 $Y=728860
X1546 1335 1293 1330 1297 2 1 MXL2HS $T=495380 799800 0 180 $X=489800 $Y=794380
X1547 1309 1275 1344 1288 2 1 MXL2HS $T=489800 819960 1 0 $X=489800 $Y=814540
X1548 1331 1299 1345 1349 2 1 MXL2HS $T=489800 870360 1 0 $X=489800 $Y=864940
X1549 1343 1251 1334 126 2 1 MXL2HS $T=496000 749400 1 180 $X=490420 $Y=749020
X1550 1356 1275 1326 1305 2 1 MXL2HS $T=497240 830040 0 180 $X=491660 $Y=824620
X1551 1359 1251 1352 1278 2 1 MXL2HS $T=500340 759480 0 180 $X=494760 $Y=754060
X1552 1349 1287 1363 1356 2 1 MXL2HS $T=495380 840120 0 0 $X=495380 $Y=839740
X1553 1236 1293 1347 1384 2 1 MXL2HS $T=497860 809880 1 0 $X=497860 $Y=804460
X1554 1364 1275 1373 1385 2 1 MXL2HS $T=497860 830040 1 0 $X=497860 $Y=824620
X1555 1365 1299 1355 1379 2 1 MXL2HS $T=497860 870360 1 0 $X=497860 $Y=864940
X1556 1388 1381 1353 1327 2 1 MXL2HS $T=504060 890520 0 180 $X=498480 $Y=885100
X1557 143 1299 1328 1351 2 1 MXL2HS $T=504680 890520 1 180 $X=499100 $Y=890140
X1558 1379 1287 1394 1364 2 1 MXL2HS $T=500960 850200 0 0 $X=500960 $Y=849820
X1559 1393 1346 1386 141 2 1 MXL2HS $T=507160 729240 1 180 $X=501580 $Y=728860
X1560 1401 1396 1387 138 2 1 MXL2HS $T=508400 769560 1 180 $X=502820 $Y=769180
X1561 1385 1293 1402 1401 2 1 MXL2HS $T=504680 809880 1 0 $X=504680 $Y=804460
X1562 1406 1381 145 1307 2 1 MXL2HS $T=510260 900600 0 180 $X=504680 $Y=895180
X1563 1384 1293 1404 148 2 1 MXL2HS $T=505300 799800 0 0 $X=505300 $Y=799420
X1564 1412 146 1390 144 2 1 MXL2HS $T=511500 739320 1 180 $X=505920 $Y=738940
X1565 1418 1381 1400 1388 2 1 MXL2HS $T=512740 890520 0 180 $X=507160 $Y=885100
X1566 1413 1396 1407 1393 2 1 MXL2HS $T=513360 769560 0 180 $X=507780 $Y=764140
X1567 1421 1416 1350 1365 2 1 MXL2HS $T=513360 870360 1 180 $X=507780 $Y=869980
X1568 1426 1419 1391 147 2 1 MXL2HS $T=513980 759480 0 180 $X=508400 $Y=754060
X1569 1409 1282 1420 1417 2 1 MXL2HS $T=516460 819960 0 180 $X=510880 $Y=814540
X1570 1417 1282 1430 1426 2 1 MXL2HS $T=511500 799800 0 0 $X=511500 $Y=799420
X1571 1432 1436 1405 1423 2 1 MXL2HS $T=517080 840120 1 180 $X=511500 $Y=839740
X1572 1423 1436 1410 1409 2 1 MXL2HS $T=518940 830040 1 180 $X=513360 $Y=829660
X1573 1448 1436 1411 1432 2 1 MXL2HS $T=518940 850200 1 180 $X=513360 $Y=849820
X1574 157 146 1440 151 2 1 MXL2HS $T=519560 719160 1 180 $X=513980 $Y=718780
X1575 1450 1416 1442 1421 2 1 MXL2HS $T=519560 880440 0 180 $X=513980 $Y=875020
X1576 1452 1381 154 1406 2 1 MXL2HS $T=519560 900600 0 180 $X=513980 $Y=895180
X1577 1437 146 1445 158 2 1 MXL2HS $T=514600 729240 0 0 $X=514600 $Y=728860
X1578 1438 1419 1446 159 2 1 MXL2HS $T=514600 749400 0 0 $X=514600 $Y=749020
X1579 1314 1444 1424 160 2 1 MXL2HS $T=515840 779640 0 0 $X=515840 $Y=779260
X1580 155 1416 1456 1464 2 1 MXL2HS $T=517700 870360 0 0 $X=517700 $Y=869980
X1581 1455 1419 1461 150 2 1 MXL2HS $T=525140 749400 0 180 $X=519560 $Y=743980
X1582 1476 1419 1462 1437 2 1 MXL2HS $T=526380 749400 1 180 $X=520800 $Y=749020
X1583 1480 1459 1467 1418 2 1 MXL2HS $T=526380 890520 0 180 $X=520800 $Y=885100
X1584 1477 1282 1441 1463 2 1 MXL2HS $T=527000 799800 1 180 $X=521420 $Y=799420
X1585 1485 1444 1433 1438 2 1 MXL2HS $T=527620 779640 1 180 $X=522040 $Y=779260
X1586 1488 1459 1475 1450 2 1 MXL2HS $T=528240 880440 1 180 $X=522660 $Y=880060
X1587 1470 163 1486 161 2 1 MXL2HS $T=523900 729240 0 0 $X=523900 $Y=728860
X1588 1479 1483 1482 1477 2 1 MXL2HS $T=529480 819960 0 180 $X=523900 $Y=814540
X1589 1494 1490 1472 1448 2 1 MXL2HS $T=529480 860280 1 180 $X=523900 $Y=859900
X1590 1464 1483 1425 1497 2 1 MXL2HS $T=524520 830040 1 0 $X=524520 $Y=824620
X1591 1498 1436 1465 1479 2 1 MXL2HS $T=530100 840120 0 180 $X=524520 $Y=834700
X1592 1463 1444 1471 1485 2 1 MXL2HS $T=525140 789720 0 0 $X=525140 $Y=789340
X1593 1502 1459 1484 1452 2 1 MXL2HS $T=531340 890520 1 180 $X=525760 $Y=890140
X1594 1510 1444 1495 164 2 1 MXL2HS $T=533200 769560 1 180 $X=527620 $Y=769180
X1595 1514 1490 1474 1499 2 1 MXL2HS $T=533820 850200 0 180 $X=528240 $Y=844780
X1596 1520 1483 1511 1503 2 1 MXL2HS $T=536300 809880 1 180 $X=530720 $Y=809500
X1597 1526 1444 1491 1510 2 1 MXL2HS $T=536920 779640 1 180 $X=531340 $Y=779260
X1598 1503 1444 1519 1526 2 1 MXL2HS $T=531340 789720 0 0 $X=531340 $Y=789340
X1599 1499 1483 1523 1520 2 1 MXL2HS $T=531960 819960 0 0 $X=531960 $Y=819580
X1600 1530 1490 1505 1494 2 1 MXL2HS $T=538780 860280 1 180 $X=533200 $Y=859900
X1601 1546 1512 1516 1498 2 1 MXL2HS $T=541260 840120 0 180 $X=535680 $Y=834700
X1602 1547 1459 170 1502 2 1 MXL2HS $T=541260 890520 1 180 $X=535680 $Y=890140
X1603 169 1490 1545 1539 2 1 MXL2HS $T=536920 870360 1 0 $X=536920 $Y=864940
X1604 1528 1551 1501 167 2 1 MXL2HS $T=543120 759480 0 180 $X=537540 $Y=754060
X1605 1539 1512 1524 1550 2 1 MXL2HS $T=538160 840120 0 0 $X=538160 $Y=839740
X1606 1567 1562 1554 1549 2 1 MXL2HS $T=545600 799800 1 180 $X=540020 $Y=799420
X1607 1550 1541 1563 1567 2 1 MXL2HS $T=540020 809880 0 0 $X=540020 $Y=809500
X1608 173 163 1556 1470 2 1 MXL2HS $T=546840 729240 0 180 $X=541260 $Y=723820
X1609 1574 1459 1560 1480 2 1 MXL2HS $T=546840 890520 0 180 $X=541260 $Y=885100
X1610 1577 1551 1558 1359 2 1 MXL2HS $T=547460 759480 1 180 $X=541880 $Y=759100
X1611 1582 1490 1564 1514 2 1 MXL2HS $T=548080 850200 1 180 $X=542500 $Y=849820
X1612 1536 1551 1575 1584 2 1 MXL2HS $T=543120 769560 1 0 $X=543120 $Y=764140
X1613 1566 1579 1544 1536 2 1 MXL2HS $T=548700 779640 1 180 $X=543120 $Y=779260
X1614 1585 1490 1570 1530 2 1 MXL2HS $T=548700 860280 1 180 $X=543120 $Y=859900
X1615 1586 1562 1571 1566 2 1 MXL2HS $T=549320 799800 0 180 $X=543740 $Y=794380
X1616 1587 1561 1569 1343 2 1 MXL2HS $T=549940 749400 0 180 $X=544360 $Y=743980
X1617 1593 172 1583 1488 2 1 MXL2HS $T=551800 880440 0 180 $X=546220 $Y=875020
X1618 1497 1562 1576 1598 2 1 MXL2HS $T=548080 819960 1 0 $X=548080 $Y=814540
X1619 1599 1512 1572 1546 2 1 MXL2HS $T=553660 840120 0 180 $X=548080 $Y=834700
X1620 1549 1579 1596 1543 2 1 MXL2HS $T=555520 779640 1 180 $X=549940 $Y=779260
X1621 1604 172 1597 1574 2 1 MXL2HS $T=555520 890520 0 180 $X=549940 $Y=885100
X1622 1610 1606 1600 1582 2 1 MXL2HS $T=556760 850200 1 180 $X=551180 $Y=849820
X1623 1598 1562 1613 1624 2 1 MXL2HS $T=553040 809880 0 0 $X=553040 $Y=809500
X1624 1543 1579 1618 1627 2 1 MXL2HS $T=553660 769560 1 0 $X=553660 $Y=764140
X1625 1628 1622 1580 1585 2 1 MXL2HS $T=559240 860280 1 180 $X=553660 $Y=859900
X1626 1637 172 1623 1593 2 1 MXL2HS $T=561100 880440 0 180 $X=555520 $Y=875020
X1627 1638 1606 1621 1610 2 1 MXL2HS $T=561720 840120 1 180 $X=556140 $Y=839740
X1628 1640 1561 1617 1535 2 1 MXL2HS $T=562340 739320 0 180 $X=556760 $Y=733900
X1629 1584 1561 1620 1641 2 1 MXL2HS $T=556760 749400 0 0 $X=556760 $Y=749020
X1630 1644 172 1633 1547 2 1 MXL2HS $T=562960 900600 0 180 $X=557380 $Y=895180
X1631 1594 1562 1629 1639 2 1 MXL2HS $T=558000 799800 0 0 $X=558000 $Y=799420
X1632 1641 1647 1619 178 2 1 MXL2HS $T=565440 729240 0 180 $X=559860 $Y=723820
X1633 1639 1579 1643 1529 2 1 MXL2HS $T=565440 779640 1 180 $X=559860 $Y=779260
X1634 1651 1606 1626 1599 2 1 MXL2HS $T=565440 830040 1 180 $X=559860 $Y=829660
X1635 1529 1579 1648 1654 2 1 MXL2HS $T=560480 769560 1 0 $X=560480 $Y=764140
X1636 1656 1561 1642 1313 2 1 MXL2HS $T=566680 739320 1 180 $X=561100 $Y=738940
X1637 1662 1562 1650 1586 2 1 MXL2HS $T=567920 799800 0 180 $X=562340 $Y=794380
X1638 1664 1622 1652 1628 2 1 MXL2HS $T=568540 860280 0 180 $X=562960 $Y=854860
X1639 1627 1659 1671 1679 2 1 MXL2HS $T=565440 749400 0 0 $X=565440 $Y=749020
X1640 1684 1606 1667 1638 2 1 MXL2HS $T=571640 840120 1 180 $X=566060 $Y=839740
X1641 1624 1669 1649 1691 2 1 MXL2HS $T=567300 779640 0 0 $X=567300 $Y=779260
X1642 1654 1659 1688 1658 2 1 MXL2HS $T=569160 759480 0 0 $X=569160 $Y=759100
X1643 1701 1661 1690 1664 2 1 MXL2HS $T=575360 860280 0 180 $X=569780 $Y=854860
X1644 1702 1661 1694 1657 2 1 MXL2HS $T=575980 860280 1 180 $X=570400 $Y=859900
X1645 1708 1659 1697 1577 2 1 MXL2HS $T=577220 749400 1 180 $X=571640 $Y=749020
X1646 1711 1647 1686 1656 2 1 MXL2HS $T=577840 729240 1 180 $X=572260 $Y=728860
X1647 1712 1669 1689 1528 2 1 MXL2HS $T=577840 779640 0 180 $X=572260 $Y=774220
X1648 1713 1710 1699 1662 2 1 MXL2HS $T=578460 799800 0 180 $X=572880 $Y=794380
X1649 1714 1710 1673 1329 2 1 MXL2HS $T=578460 809880 1 180 $X=572880 $Y=809500
X1650 1719 1710 1705 1300 2 1 MXL2HS $T=579700 809880 0 180 $X=574120 $Y=804460
X1651 1721 184 1707 1644 2 1 MXL2HS $T=579700 900600 0 180 $X=574120 $Y=895180
X1652 1729 1669 1704 1413 2 1 MXL2HS $T=581560 779640 1 180 $X=575980 $Y=779260
X1653 1732 1728 1715 1692 2 1 MXL2HS $T=582180 870360 1 180 $X=576600 $Y=869980
X1654 1679 1647 1730 1738 2 1 MXL2HS $T=577840 729240 0 0 $X=577840 $Y=728860
X1655 1747 1710 1727 1713 2 1 MXL2HS $T=585280 799800 0 180 $X=579700 $Y=794380
X1656 189 1647 1740 1565 2 1 MXL2HS $T=586520 719160 1 180 $X=580940 $Y=718780
X1657 1754 1710 1743 1594 2 1 MXL2HS $T=587760 809880 1 180 $X=582180 $Y=809500
X1658 1755 1728 1736 1721 2 1 MXL2HS $T=587760 880440 1 180 $X=582180 $Y=880060
X1659 191 1745 1748 1708 2 1 MXL2HS $T=588380 729240 0 180 $X=582800 $Y=723820
X1660 1761 1669 1749 1455 2 1 MXL2HS $T=589000 769560 1 180 $X=583420 $Y=769180
X1661 1765 1669 1752 1476 2 1 MXL2HS $T=589620 779640 0 180 $X=584040 $Y=774220
X1662 1658 1659 1759 1766 2 1 MXL2HS $T=584660 749400 0 0 $X=584660 $Y=749020
X1663 1691 1659 1734 1767 2 1 MXL2HS $T=584660 759480 1 0 $X=584660 $Y=754060
X1664 1773 1728 1718 1732 2 1 MXL2HS $T=592100 870360 0 180 $X=586520 $Y=864940
X1665 1779 1776 1744 1731 2 1 MXL2HS $T=593340 830040 0 180 $X=587760 $Y=824620
X1666 1788 1710 1760 1747 2 1 MXL2HS $T=597060 799800 0 180 $X=591480 $Y=794380
X1667 1789 1728 1780 1755 2 1 MXL2HS $T=597060 870360 1 180 $X=591480 $Y=869980
X1668 1767 1745 1769 1794 2 1 MXL2HS $T=592100 749400 0 0 $X=592100 $Y=749020
X1669 1795 1790 1784 1335 2 1 MXL2HS $T=598300 799800 1 180 $X=592720 $Y=799420
X1670 1766 1745 1778 1797 2 1 MXL2HS $T=593340 749400 1 0 $X=593340 $Y=743980
X1671 1801 1796 1787 1702 2 1 MXL2HS $T=599540 860280 1 180 $X=593960 $Y=859900
X1672 1804 194 1783 197 2 1 MXL2HS $T=600780 890520 1 180 $X=595200 $Y=890140
X1673 1812 1776 1791 1779 2 1 MXL2HS $T=601400 830040 0 180 $X=595820 $Y=824620
X1674 1808 1790 1802 1788 2 1 MXL2HS $T=602640 789720 1 180 $X=597060 $Y=789340
X1675 1824 1790 1814 1808 2 1 MXL2HS $T=604500 789720 0 180 $X=598920 $Y=784300
X1676 1831 1796 1817 1789 2 1 MXL2HS $T=605740 870360 0 180 $X=600160 $Y=864940
X1677 1832 1826 1818 1804 2 1 MXL2HS $T=605740 880440 1 180 $X=600160 $Y=880060
X1678 1836 1827 1792 1735 2 1 MXL2HS $T=606360 840120 0 180 $X=600780 $Y=834700
X1679 1797 1833 1822 1819 2 1 MXL2HS $T=606980 749400 1 180 $X=601400 $Y=749020
X1680 1841 1776 1810 1823 2 1 MXL2HS $T=607600 819960 1 180 $X=602020 $Y=819580
X1681 1823 194 1834 203 2 1 MXL2HS $T=602020 890520 0 0 $X=602020 $Y=890140
X1682 1738 1745 1799 1847 2 1 MXL2HS $T=603260 739320 1 0 $X=603260 $Y=733900
X1683 1819 1790 1851 1824 2 1 MXL2HS $T=605740 769560 0 0 $X=605740 $Y=769180
X1684 1846 1796 1858 1801 2 1 MXL2HS $T=606360 860280 1 0 $X=606360 $Y=854860
X1685 1870 1827 1856 1812 2 1 MXL2HS $T=613800 830040 0 180 $X=608220 $Y=824620
X1686 1855 1868 1859 1841 2 1 MXL2HS $T=614420 809880 0 180 $X=608840 $Y=804460
X1687 1865 1826 1853 205 2 1 MXL2HS $T=614420 900600 0 180 $X=608840 $Y=895180
X1688 208 1745 1839 1711 2 1 MXL2HS $T=615040 729240 1 180 $X=609460 $Y=728860
X1689 1847 1833 1825 1862 2 1 MXL2HS $T=615660 749400 1 180 $X=610080 $Y=749020
X1690 1876 1827 1857 1836 2 1 MXL2HS $T=616280 840120 0 180 $X=610700 $Y=834700
X1691 1878 1776 1872 1865 2 1 MXL2HS $T=616900 819960 1 180 $X=611320 $Y=819580
X1692 1879 1827 1869 1803 2 1 MXL2HS $T=616900 850200 0 180 $X=611320 $Y=844780
X1693 1862 1790 1871 1887 2 1 MXL2HS $T=613180 769560 1 0 $X=613180 $Y=764140
X1694 1873 1868 1881 1892 2 1 MXL2HS $T=614420 799800 0 0 $X=614420 $Y=799420
X1695 1880 1826 1864 211 2 1 MXL2HS $T=615040 870360 0 0 $X=615040 $Y=869980
X1696 1892 1868 1884 1880 2 1 MXL2HS $T=621240 819960 0 180 $X=615660 $Y=814540
X1697 214 1899 1867 1873 2 1 MXL2HS $T=623100 729240 0 180 $X=617520 $Y=723820
X1698 1913 1883 1852 1855 2 1 MXL2HS $T=624340 779640 1 180 $X=618760 $Y=779260
X1699 1914 1909 1901 1832 2 1 MXL2HS $T=624340 880440 0 180 $X=618760 $Y=875020
X1700 212 1899 1889 1895 2 1 MXL2HS $T=619380 739320 1 0 $X=619380 $Y=733900
X1701 1794 1833 1910 1885 2 1 MXL2HS $T=620000 749400 0 0 $X=620000 $Y=749020
X1702 1897 1826 1915 218 2 1 MXL2HS $T=620000 880440 0 0 $X=620000 $Y=880060
X1703 1895 1868 1874 1878 2 1 MXL2HS $T=626200 799800 1 180 $X=620620 $Y=799420
X1704 1923 1917 1904 1897 2 1 MXL2HS $T=626200 809880 0 180 $X=620620 $Y=804460
X1705 1929 1921 1911 1830 2 1 MXL2HS $T=626820 850200 0 180 $X=621240 $Y=844780
X1706 1930 1920 1912 1831 2 1 MXL2HS $T=626820 860280 1 180 $X=621240 $Y=859900
X1707 1933 1883 1926 1923 2 1 MXL2HS $T=630540 769560 1 180 $X=624960 $Y=769180
X1708 1941 1921 1931 1928 2 1 MXL2HS $T=630540 840120 0 180 $X=624960 $Y=834700
X1709 222 1899 1925 1933 2 1 MXL2HS $T=631780 729240 0 180 $X=626200 $Y=723820
X1710 1885 1932 1944 1913 2 1 MXL2HS $T=626820 759480 0 0 $X=626820 $Y=759100
X1711 1928 219 1918 221 2 1 MXL2HS $T=632400 900600 0 180 $X=626820 $Y=895180
X1712 1954 1920 1922 1846 2 1 MXL2HS $T=633640 860280 1 180 $X=628060 $Y=859900
X1713 226 1899 1948 1945 2 1 MXL2HS $T=634880 739320 0 180 $X=629300 $Y=733900
X1714 1945 1955 1946 1941 2 1 MXL2HS $T=634880 809880 0 180 $X=629300 $Y=804460
X1715 1887 1955 1939 1950 2 1 MXL2HS $T=636740 789720 1 180 $X=631160 $Y=789340
X1716 224 1932 1949 1970 2 1 MXL2HS $T=632400 759480 0 0 $X=632400 $Y=759100
X1717 232 219 227 1754 2 1 MXL2HS $T=639220 900600 0 180 $X=633640 $Y=895180
X1718 1976 1917 1958 1961 2 1 MXL2HS $T=639840 819960 0 180 $X=634260 $Y=814540
X1719 1964 1955 1974 1985 2 1 MXL2HS $T=634880 799800 0 0 $X=634880 $Y=799420
X1720 1989 1883 1953 1964 2 1 MXL2HS $T=641700 769560 1 180 $X=636120 $Y=769180
X1721 1961 1920 1957 229 2 1 MXL2HS $T=641700 860280 1 180 $X=636120 $Y=859900
X1722 1994 1883 1978 1976 2 1 MXL2HS $T=642940 779640 1 180 $X=637360 $Y=779260
X1723 1995 1921 1981 1876 2 1 MXL2HS $T=642940 840120 0 180 $X=637360 $Y=834700
X1724 233 230 1971 1996 2 1 MXL2HS $T=637980 729240 1 0 $X=637980 $Y=723820
X1725 1950 1917 1966 1992 2 1 MXL2HS $T=637980 830040 1 0 $X=637980 $Y=824620
X1726 1985 1920 1983 238 2 1 MXL2HS $T=639220 870360 0 0 $X=639220 $Y=869980
X1727 235 230 237 2004 2 1 MXL2HS $T=639840 719160 0 0 $X=639840 $Y=718780
X1728 2005 1955 1972 1990 2 1 MXL2HS $T=645420 799800 0 180 $X=639840 $Y=794380
X1729 1992 1921 1940 2001 2 1 MXL2HS $T=640460 850200 1 0 $X=640460 $Y=844780
X1730 2009 1999 1975 216 2 1 MXL2HS $T=646040 890520 0 180 $X=640460 $Y=885100
X1731 236 2006 1937 1989 2 1 MXL2HS $T=646660 749400 0 180 $X=641080 $Y=743980
X1732 1996 1932 1998 2014 2 1 MXL2HS $T=641700 759480 0 0 $X=641700 $Y=759100
X1733 2016 1999 2007 239 2 1 MXL2HS $T=648520 890520 1 180 $X=642940 $Y=890140
X1734 2001 1999 240 242 2 1 MXL2HS $T=642940 900600 1 0 $X=642940 $Y=895180
X1735 2023 2000 2010 1870 2 1 MXL2HS $T=650380 830040 0 180 $X=644800 $Y=824620
X1736 2008 1920 2020 243 2 1 MXL2HS $T=645420 870360 0 0 $X=645420 $Y=869980
X1737 2029 1921 2017 1879 2 1 MXL2HS $T=651620 840120 1 180 $X=646040 $Y=839740
X1738 241 2006 2024 1994 2 1 MXL2HS $T=646660 749400 1 0 $X=646660 $Y=743980
X1739 2035 1920 2015 1954 2 1 MXL2HS $T=652240 860280 0 180 $X=646660 $Y=854860
X1740 1970 1932 2033 2040 2 1 MXL2HS $T=647900 769560 1 0 $X=647900 $Y=764140
X1741 2014 1955 2013 2042 2 1 MXL2HS $T=648520 789720 0 0 $X=648520 $Y=789340
X1742 244 2006 247 2048 2 1 MXL2HS $T=650380 719160 0 0 $X=650380 $Y=718780
X1743 2051 2043 2041 1914 2 1 MXL2HS $T=656580 870360 1 180 $X=651000 $Y=869980
X1744 2004 2045 2025 2057 2 1 MXL2HS $T=652860 749400 1 0 $X=652860 $Y=743980
X1745 248 2006 2031 2005 2 1 MXL2HS $T=659060 739320 0 180 $X=653480 $Y=733900
X1746 2042 2000 2060 2064 2 1 MXL2HS $T=654720 819960 1 0 $X=654720 $Y=814540
X1747 2066 2043 2055 2016 2 1 MXL2HS $T=660920 860280 0 180 $X=655340 $Y=854860
X1748 2079 2075 2059 1930 2 1 MXL2HS $T=663400 830040 0 180 $X=657820 $Y=824620
X1749 2040 1955 2062 2080 2 1 MXL2HS $T=658440 789720 0 0 $X=658440 $Y=789340
X1750 250 2006 251 2089 2 1 MXL2HS $T=660300 719160 0 0 $X=660300 $Y=718780
X1751 2048 2045 2038 2076 2 1 MXL2HS $T=666500 749400 0 180 $X=660920 $Y=743980
X1752 2076 2049 2074 2094 2 1 MXL2HS $T=660920 769560 0 0 $X=660920 $Y=769180
X1753 2077 2000 2067 2095 2 1 MXL2HS $T=660920 819960 1 0 $X=660920 $Y=814540
X1754 2080 2043 2068 2097 2 1 MXL2HS $T=661540 850200 0 0 $X=661540 $Y=849820
X1755 2064 2083 2071 255 2 1 MXL2HS $T=662160 880440 0 0 $X=662160 $Y=880060
X1756 2057 2049 2069 2077 2 1 MXL2HS $T=663400 779640 1 0 $X=663400 $Y=774220
X1757 2112 2075 2100 2023 2 1 MXL2HS $T=670840 830040 0 180 $X=665260 $Y=824620
X1758 257 2045 2117 2110 2 1 MXL2HS $T=667740 739320 1 0 $X=667740 $Y=733900
X1759 2089 2045 2082 2124 2 1 MXL2HS $T=667740 749400 1 0 $X=667740 $Y=743980
X1760 2126 2075 2102 1995 2 1 MXL2HS $T=673320 809880 1 180 $X=667740 $Y=809500
X1761 2095 2043 2046 258 2 1 MXL2HS $T=668360 870360 1 0 $X=668360 $Y=864940
X1762 2110 2107 2120 2132 2 1 MXL2HS $T=668980 759480 0 0 $X=668980 $Y=759100
X1763 2094 2075 2114 2115 2 1 MXL2HS $T=675180 799800 1 180 $X=669600 $Y=799420
X1764 2097 2083 2056 263 2 1 MXL2HS $T=670220 890520 1 0 $X=670220 $Y=885100
X1765 2132 2135 2113 2119 2 1 MXL2HS $T=676420 779640 0 180 $X=670840 $Y=774220
X1766 2115 2123 2133 264 2 1 MXL2HS $T=670840 860280 1 0 $X=670840 $Y=854860
X1767 2119 2075 2121 2125 2 1 MXL2HS $T=677040 799800 0 180 $X=671460 $Y=794380
X1768 2125 2129 2070 2139 2 1 MXL2HS $T=671460 840120 0 0 $X=671460 $Y=839740
X1769 261 262 2137 2143 2 1 MXL2HS $T=672080 719160 0 0 $X=672080 $Y=718780
X1770 2144 2129 2131 259 2 1 MXL2HS $T=677660 830040 1 180 $X=672080 $Y=829660
X1771 2150 2123 2138 2009 2 1 MXL2HS $T=679520 860280 1 180 $X=673940 $Y=859900
X1772 2155 2135 2118 2141 2 1 MXL2HS $T=680760 779640 1 180 $X=675180 $Y=779260
X1773 265 2045 2152 2158 2 1 MXL2HS $T=675800 739320 1 0 $X=675800 $Y=733900
X1774 2124 2135 2151 2155 2 1 MXL2HS $T=675800 759480 0 0 $X=675800 $Y=759100
X1775 2161 2153 2122 2126 2 1 MXL2HS $T=682000 799800 1 180 $X=676420 $Y=799420
X1776 2141 2129 2154 2164 2 1 MXL2HS $T=677660 840120 0 0 $X=677660 $Y=839740
X1777 2139 2083 2160 2168 2 1 MXL2HS $T=677660 890520 1 0 $X=677660 $Y=885100
X1778 2175 2123 2157 267 2 1 MXL2HS $T=684480 860280 0 180 $X=678900 $Y=854860
X1779 2177 2075 2165 1929 2 1 MXL2HS $T=685720 819960 0 180 $X=680140 $Y=814540
X1780 2178 2123 2166 269 2 1 MXL2HS $T=685720 860280 1 180 $X=680140 $Y=859900
X1781 2164 2083 2145 2181 2 1 MXL2HS $T=680760 880440 0 0 $X=680760 $Y=880060
X1782 2183 274 2174 272 2 1 MXL2HS $T=686960 900600 0 180 $X=681380 $Y=895180
X1783 2185 2135 2169 2170 2 1 MXL2HS $T=687580 779640 0 180 $X=682000 $Y=774220
X1784 2170 2135 2179 2180 2 1 MXL2HS $T=682000 779640 0 0 $X=682000 $Y=779260
X1785 2186 2153 2134 2066 2 1 MXL2HS $T=688200 799800 1 180 $X=682620 $Y=799420
X1786 273 2107 2184 2193 2 1 MXL2HS $T=683240 759480 1 0 $X=683240 $Y=754060
X1787 2180 2129 2159 2196 2 1 MXL2HS $T=684480 840120 0 0 $X=684480 $Y=839740
X1788 271 2045 2194 2185 2 1 MXL2HS $T=685100 749400 1 0 $X=685100 $Y=743980
X1789 2196 2083 2198 2210 2 1 MXL2HS $T=688200 880440 1 0 $X=688200 $Y=875020
X1790 2214 2209 2197 2079 2 1 MXL2HS $T=694400 809880 1 180 $X=688820 $Y=809500
X1791 2220 2209 2190 2047 2 1 MXL2HS $T=696260 799800 1 180 $X=690680 $Y=799420
X1792 2224 2129 2205 252 2 1 MXL2HS $T=697500 840120 0 180 $X=691920 $Y=834700
X1793 2230 2153 2218 1729 2 1 MXL2HS $T=699360 789720 1 180 $X=693780 $Y=789340
X1794 2231 2227 2207 2178 2 1 MXL2HS $T=699360 850200 1 180 $X=693780 $Y=849820
X1795 2168 2208 2173 2240 2 1 MXL2HS $T=696260 890520 1 0 $X=696260 $Y=885100
X1796 2181 2208 2187 2251 2 1 MXL2HS $T=698120 880440 0 0 $X=698120 $Y=880060
X1797 2264 2227 2254 2175 2 1 MXL2HS $T=706800 840120 0 180 $X=701220 $Y=834700
X1798 2269 2267 2260 2224 2 1 MXL2HS $T=709280 819960 1 180 $X=703700 $Y=819580
X1799 2273 2267 2266 1795 2 1 MXL2HS $T=710520 809880 1 180 $X=704940 $Y=809500
X1800 2278 2227 2245 2035 2 1 MXL2HS $T=711140 860280 0 180 $X=705560 $Y=854860
X1801 2210 2208 2272 2281 2 1 MXL2HS $T=706180 880440 0 0 $X=706180 $Y=880060
X1802 2292 2209 2274 1712 2 1 MXL2HS $T=713620 789720 1 180 $X=708040 $Y=789340
X1803 2240 2275 2286 2295 2 1 MXL2HS $T=708660 890520 1 0 $X=708660 $Y=885100
X1804 2299 2267 2284 2177 2 1 MXL2HS $T=714860 809880 0 180 $X=709280 $Y=804460
X1805 2306 2267 2270 2112 2 1 MXL2HS $T=716100 819960 1 180 $X=710520 $Y=819580
X1806 2307 2300 2291 2183 2 1 MXL2HS $T=716100 870360 0 180 $X=710520 $Y=864940
X1807 2251 2208 2285 300 2 1 MXL2HS $T=711760 880440 0 0 $X=711760 $Y=880060
X1808 2308 2300 2237 2051 2 1 MXL2HS $T=717960 870360 1 180 $X=712380 $Y=869980
X1809 2281 2275 2317 307 2 1 MXL2HS $T=719200 890520 0 0 $X=719200 $Y=890140
X1810 2316 2319 2333 2323 2 1 MXL2HS $T=725400 749400 1 180 $X=719820 $Y=749020
X1811 2348 2320 2337 2294 2 1 MXL2HS $T=726020 850200 0 180 $X=720440 $Y=844780
X1812 2350 2320 2342 2144 2 1 MXL2HS $T=726640 830040 1 180 $X=721060 $Y=829660
X1813 2351 2300 2343 2308 2 1 MXL2HS $T=726640 870360 1 180 $X=721060 $Y=869980
X1814 2345 2320 2341 2150 2 1 MXL2HS $T=728500 830040 0 180 $X=722920 $Y=824620
X1815 2359 2320 2322 2231 2 1 MXL2HS $T=729120 850200 1 180 $X=723540 $Y=849820
X1816 2363 2300 2353 2268 2 1 MXL2HS $T=730360 860280 1 180 $X=724780 $Y=859900
X1817 2379 2378 2369 2306 2 1 MXL2HS $T=734080 830040 1 180 $X=728500 $Y=829660
X1818 2399 2320 2376 2278 2 1 MXL2HS $T=738420 850200 1 180 $X=732840 $Y=849820
X1819 2405 2378 2394 2292 2 1 MXL2HS $T=739660 830040 0 180 $X=734080 $Y=824620
X1820 2295 2275 2398 328 2 1 MXL2HS $T=734080 890520 0 0 $X=734080 $Y=890140
X1821 2426 2378 2404 2230 2 1 MXL2HS $T=744620 799800 1 180 $X=739040 $Y=799420
X1822 2436 2430 2418 2345 2 1 MXL2HS $T=746480 830040 0 180 $X=740900 $Y=824620
X1823 2444 2430 2421 2264 2 1 MXL2HS $T=748340 840120 0 180 $X=742760 $Y=834700
X1824 2438 2300 2453 2463 2 1 MXL2HS $T=745240 880440 0 0 $X=745240 $Y=880060
X1825 2464 2430 2431 2444 2 1 MXL2HS $T=752060 850200 1 180 $X=746480 $Y=849820
X1826 340 2300 2448 2438 2 1 MXL2HS $T=753300 890520 1 180 $X=747720 $Y=890140
X1827 2483 2378 2455 2299 2 1 MXL2HS $T=755780 809880 1 180 $X=750200 $Y=809500
X1828 2491 2430 2475 2379 2 1 MXL2HS $T=757020 840120 0 180 $X=751440 $Y=834700
X1829 2497 2430 2480 2350 2 1 MXL2HS $T=758260 830040 0 180 $X=752680 $Y=824620
X1830 2504 2474 2486 2289 2 1 MXL2HS $T=758880 799800 0 180 $X=753300 $Y=794380
X1831 2463 2430 2411 2405 2 1 MXL2HS $T=754540 850200 1 0 $X=754540 $Y=844780
X1832 2492 2508 2460 2464 2 1 MXL2HS $T=760740 880440 1 180 $X=755160 $Y=880060
X1833 2512 2508 345 2492 2 1 MXL2HS $T=760740 890520 1 180 $X=755160 $Y=890140
X1834 2525 2508 2440 2351 2 1 MXL2HS $T=763220 880440 0 180 $X=757640 $Y=875020
X1835 2530 2487 2515 2214 2 1 MXL2HS $T=763840 819960 1 180 $X=758260 $Y=819580
X1836 350 2435 2481 2491 2 1 MXL2HS $T=763840 870360 0 180 $X=758260 $Y=864940
X1837 2544 2487 2484 2161 2 1 MXL2HS $T=766940 809880 0 180 $X=761360 $Y=804460
X1838 2548 2487 2532 2269 2 1 MXL2HS $T=767560 809880 1 180 $X=761980 $Y=809500
X1839 2570 2435 2555 2399 2 1 MXL2HS $T=770660 850200 1 180 $X=765080 $Y=849820
X1840 356 2508 2534 2363 2 1 MXL2HS $T=770660 880440 1 180 $X=765080 $Y=880060
X1841 2591 2435 2575 2348 2 1 MXL2HS $T=774380 850200 0 180 $X=768800 $Y=844780
X1842 2593 2435 2566 2359 2 1 MXL2HS $T=775000 860280 0 180 $X=769420 $Y=854860
X1843 2595 2474 2552 2318 2 1 MXL2HS $T=775620 799800 1 180 $X=770040 $Y=799420
X1844 358 2508 2556 2525 2 1 MXL2HS $T=776240 890520 1 180 $X=770660 $Y=890140
X1845 2604 2553 2561 2443 2 1 MXL2HS $T=778100 809880 1 180 $X=772520 $Y=809500
X1846 2607 2553 2554 2273 2 1 MXL2HS $T=778720 830040 0 180 $X=773140 $Y=824620
X1847 2629 2474 2618 2504 2 1 MXL2HS $T=783680 799800 1 180 $X=778100 $Y=799420
X1848 362 2589 2616 2600 2 1 MXL2HS $T=783680 880440 1 180 $X=778100 $Y=880060
X1849 2634 2553 2622 2415 2 1 MXL2HS $T=784920 830040 0 180 $X=779340 $Y=824620
X1850 363 2589 2602 2570 2 1 MXL2HS $T=784920 890520 1 180 $X=779340 $Y=890140
X1851 367 2589 2598 2591 2 1 MXL2HS $T=788640 870360 0 180 $X=783060 $Y=864940
X1852 2672 2643 2642 2548 2 1 MXL2HS $T=792980 809880 0 180 $X=787400 $Y=804460
X1853 371 369 2659 2593 2 1 MXL2HS $T=793600 890520 1 180 $X=788020 $Y=890140
X1854 370 2666 2652 2634 2 1 MXL2HS $T=794220 860280 0 180 $X=788640 $Y=854860
X1855 372 2666 2655 2626 2 1 MXL2HS $T=794840 840120 1 180 $X=789260 $Y=839740
X1856 2686 2680 2676 2530 2 1 MXL2HS $T=796700 819960 1 180 $X=791120 $Y=819580
X1857 374 2666 2653 2629 2 1 MXL2HS $T=797940 870360 1 180 $X=792360 $Y=869980
X1858 2708 2643 2697 2544 2 1 MXL2HS $T=801660 809880 1 180 $X=796080 $Y=809500
X1859 2711 2680 2701 2497 2 1 MXL2HS $T=802280 830040 0 180 $X=796700 $Y=824620
X1860 377 2666 2702 2694 2 1 MXL2HS $T=802280 850200 1 180 $X=796700 $Y=849820
X1861 384 2680 2714 2672 2 1 MXL2HS $T=806000 840120 1 180 $X=800420 $Y=839740
X1862 2705 2643 2718 2595 2 1 MXL2HS $T=806620 809880 0 180 $X=801040 $Y=804460
X1863 379 369 383 384 2 1 MXL2HS $T=801040 900600 1 0 $X=801040 $Y=895180
X1864 387 2716 2733 2708 2 1 MXL2HS $T=809100 870360 1 180 $X=803520 $Y=869980
X1865 390 2716 2739 2711 2 1 MXL2HS $T=811580 880440 1 180 $X=806000 $Y=880060
X1866 401 2811 2819 2828 2 1 MXL2HS $T=823360 779640 0 0 $X=823360 $Y=779260
X1867 281 2811 2773 2829 2 1 MXL2HS $T=823980 799800 1 0 $X=823980 $Y=794380
X1868 405 2811 2802 2845 2 1 MXL2HS $T=825840 779640 1 0 $X=825840 $Y=774220
X1869 2829 2832 2807 2859 2 1 MXL2HS $T=827080 819960 0 0 $X=827080 $Y=819580
X1870 2828 2832 2822 2865 2 1 MXL2HS $T=828940 809880 1 0 $X=828940 $Y=804460
X1871 2193 2811 2877 2883 2 1 MXL2HS $T=833280 799800 1 0 $X=833280 $Y=794380
X1872 415 2811 2874 2894 2 1 MXL2HS $T=836380 779640 1 0 $X=836380 $Y=774220
X1873 2845 2832 2878 2908 2 1 MXL2HS $T=839480 809880 0 0 $X=839480 $Y=809500
X1874 2894 2832 2919 2954 2 1 MXL2HS $T=847540 809880 1 0 $X=847540 $Y=804460
X1875 2883 2832 2945 2955 2 1 MXL2HS $T=847540 819960 1 0 $X=847540 $Y=814540
X1876 2143 3003 3013 3024 2 1 MXL2HS $T=859320 799800 0 0 $X=859320 $Y=799420
X1877 3024 3003 3016 3004 2 1 MXL2HS $T=866760 809880 0 180 $X=861180 $Y=804460
X1878 2158 3003 3031 3043 2 1 MXL2HS $T=861800 799800 1 0 $X=861800 $Y=794380
X1879 3043 3003 3055 3096 2 1 MXL2HS $T=869860 809880 0 0 $X=869860 $Y=809500
X1880 452 3003 3125 3135 2 1 MXL2HS $T=876680 809880 1 0 $X=876680 $Y=804460
X1881 3135 3003 3129 3128 2 1 MXL2HS $T=884740 809880 1 180 $X=879160 $Y=809500
X1882 3122 3133 3048 3115 2 1 MXL2HS $T=879780 789720 1 0 $X=879780 $Y=784300
X1883 3529 3528 3538 3546 2 1 MXL2HS $T=949220 880440 0 0 $X=949220 $Y=880060
X1884 104 27 1 2 INV12CK $T=461280 890520 0 180 $X=451360 $Y=885100
X1885 1338 882 1 2 INV12CK $T=491660 809880 0 0 $X=491660 $Y=809500
X1886 1338 1339 1 2 INV12CK $T=561100 809880 0 0 $X=561100 $Y=809500
X1887 201 1733 1 2 INV12CK $T=599540 729240 0 0 $X=599540 $Y=728860
X1888 104 198 1 2 INV12CK $T=616280 890520 0 180 $X=606360 $Y=885100
X1889 215 210 1 2 INV12CK $T=623100 759480 1 180 $X=613180 $Y=759100
X1890 1942 104 1 2 INV12CK $T=629920 890520 0 180 $X=620000 $Y=885100
X1891 1942 1338 1 2 INV12CK $T=655340 809880 0 0 $X=655340 $Y=809500
X1892 249 1942 1 2 INV12CK $T=657820 799800 0 0 $X=657820 $Y=799420
X1893 1942 253 1 2 INV12CK $T=667740 890520 0 180 $X=657820 $Y=885100
X1894 1338 2127 1 2 INV12CK $T=678900 819960 0 180 $X=668980 $Y=814540
X1895 253 270 1 2 INV12CK $T=685100 880440 0 180 $X=675180 $Y=875020
X1896 3155 2687 1 2 INV12CK $T=886600 779640 0 180 $X=876680 $Y=774220
X1897 457 3155 1 2 INV12CK $T=881640 739320 0 0 $X=881640 $Y=738940
X1898 3155 557 1 2 INV12CK $T=982080 739320 0 0 $X=982080 $Y=738940
X1899 3155 3649 1 2 INV12CK $T=983320 759480 0 0 $X=983320 $Y=759100
X1900 612 602 1 2 604 AN2 $T=317440 749400 0 180 $X=314960 $Y=743980
X1901 645 648 1 2 651 AN2 $T=327980 739320 0 0 $X=327980 $Y=738940
X1902 680 676 1 2 653 AN2 $T=336040 809880 0 180 $X=333560 $Y=804460
X1903 936 918 1 2 905 AN2 $T=397420 759480 1 180 $X=394940 $Y=759100
X1904 1206 1157 1 2 114 AN2 $T=468720 719160 0 0 $X=468720 $Y=718780
X1905 2536 2522 1 2 2559 AN2 $T=765080 759480 0 0 $X=765080 $Y=759100
X1906 2946 2937 1 2 2922 AN2 $T=850640 860280 0 180 $X=848160 $Y=854860
X1907 2978 2974 1 2 2927 AN2 $T=856840 759480 0 180 $X=854360 $Y=754060
X1908 3198 3230 1 2 3058 AN2 $T=899620 769560 0 180 $X=897140 $Y=764140
X1909 3641 3638 1 2 554 AN2 $T=982700 719160 1 180 $X=980220 $Y=718780
X1910 592 590 594 1 2 ND2 $T=306900 759480 1 0 $X=306900 $Y=754060
X1911 597 593 600 1 2 ND2 $T=311860 739320 0 0 $X=311860 $Y=738940
X1912 629 602 632 1 2 ND2 $T=323020 759480 1 0 $X=323020 $Y=754060
X1913 637 594 641 1 2 ND2 $T=324880 759480 0 0 $X=324880 $Y=759100
X1914 631 609 646 1 2 ND2 $T=327360 769560 0 0 $X=327360 $Y=769180
X1915 652 645 656 1 2 ND2 $T=329220 749400 1 0 $X=329220 $Y=743980
X1916 654 632 658 1 2 ND2 $T=329840 759480 1 0 $X=329840 $Y=754060
X1917 664 637 659 1 2 ND2 $T=332940 759480 1 180 $X=331080 $Y=759100
X1918 663 654 671 1 2 ND2 $T=332320 759480 1 0 $X=332320 $Y=754060
X1919 673 659 668 1 2 ND2 $T=334800 759480 1 180 $X=332940 $Y=759100
X1920 684 646 677 1 2 ND2 $T=337280 779640 1 0 $X=337280 $Y=774220
X1921 688 658 682 1 2 ND2 $T=337900 759480 1 0 $X=337900 $Y=754060
X1922 705 626 709 1 2 ND2 $T=341620 799800 0 0 $X=341620 $Y=799420
X1923 708 681 712 1 2 ND2 $T=342240 779640 0 0 $X=342240 $Y=779260
X1924 714 676 706 1 2 ND2 $T=344720 809880 1 0 $X=344720 $Y=804460
X1925 694 19 698 1 2 ND2 $T=345340 729240 1 0 $X=345340 $Y=723820
X1926 720 726 722 1 2 ND2 $T=350300 759480 1 180 $X=348440 $Y=759100
X1927 726 707 733 1 2 ND2 $T=350300 759480 0 0 $X=350300 $Y=759100
X1928 734 723 730 1 2 ND2 $T=354640 799800 0 0 $X=354640 $Y=799420
X1929 820 805 775 1 2 ND2 $T=373240 789720 0 180 $X=371380 $Y=784300
X1930 850 884 837 1 2 ND2 $T=383780 789720 0 0 $X=383780 $Y=789340
X1931 881 856 864 1 2 ND2 $T=385640 729240 1 0 $X=385640 $Y=723820
X1932 884 889 878 1 2 ND2 $T=386260 789720 0 0 $X=386260 $Y=789340
X1933 942 936 950 1 2 ND2 $T=398660 759480 1 0 $X=398660 $Y=754060
X1934 976 975 892 1 2 ND2 $T=405480 769560 1 0 $X=405480 $Y=764140
X1935 976 901 982 1 2 ND2 $T=405480 769560 0 0 $X=405480 $Y=769180
X1936 965 920 53 1 2 ND2 $T=407960 759480 1 0 $X=407960 $Y=754060
X1937 70 1046 1039 1 2 ND2 $T=424080 779640 0 180 $X=422220 $Y=774220
X1938 1041 804 1067 1 2 ND2 $T=423460 769560 0 0 $X=423460 $Y=769180
X1939 1056 1067 1045 1 2 ND2 $T=424700 769560 1 0 $X=424700 $Y=764140
X1940 75 79 63 1 2 ND2 $T=432140 719160 1 180 $X=430280 $Y=718780
X1941 44 1094 1098 1 2 ND2 $T=434000 719160 0 0 $X=434000 $Y=718780
X1942 2235 2226 2195 1 2 ND2 $T=700600 729240 1 180 $X=698740 $Y=728860
X1943 2298 2311 2305 1 2 ND2 $T=713620 749400 0 0 $X=713620 $Y=749020
X1944 298 2312 2282 1 2 ND2 $T=717340 759480 0 180 $X=715480 $Y=754060
X1945 2408 2400 2327 1 2 ND2 $T=739660 739320 0 180 $X=737800 $Y=733900
X1946 2330 2410 2407 1 2 ND2 $T=744000 769560 0 0 $X=744000 $Y=769180
X1947 2535 2545 2434 1 2 ND2 $T=766320 749400 1 180 $X=764460 $Y=749020
X1948 2584 2587 2526 1 2 ND2 $T=773140 769560 0 0 $X=773140 $Y=769180
X1949 2590 378 2695 1 2 ND2 $T=799800 719160 1 180 $X=797940 $Y=718780
X1950 2679 2712 2650 1 2 ND2 $T=800420 739320 0 180 $X=798560 $Y=733900
X1951 2790 2803 2758 1 2 ND2 $T=823980 729240 1 180 $X=822120 $Y=728860
X1952 2772 2794 2799 1 2 ND2 $T=822120 860280 1 0 $X=822120 $Y=854860
X1953 2797 2769 2780 1 2 ND2 $T=823360 739320 1 0 $X=823360 $Y=733900
X1954 2781 2805 2806 1 2 ND2 $T=825220 759480 1 0 $X=825220 $Y=754060
X1955 2831 2844 2834 1 2 ND2 $T=831420 749400 1 0 $X=831420 $Y=743980
X1956 2827 2834 2817 1 2 ND2 $T=832660 749400 0 0 $X=832660 $Y=749020
X1957 2881 2882 2885 1 2 ND2 $T=838240 739320 0 0 $X=838240 $Y=738940
X1958 2880 2885 2742 1 2 ND2 $T=840720 749400 1 180 $X=838860 $Y=749020
X1959 418 2901 407 1 2 ND2 $T=841960 900600 1 0 $X=841960 $Y=895180
X1960 2896 2917 2911 1 2 ND2 $T=846300 870360 1 180 $X=844440 $Y=869980
X1961 2896 2925 2915 1 2 ND2 $T=848160 880440 1 0 $X=848160 $Y=875020
X1962 2966 2967 427 1 2 ND2 $T=853740 890520 1 0 $X=853740 $Y=885100
X1963 2972 2958 433 1 2 ND2 $T=854980 860280 1 0 $X=854980 $Y=854860
X1964 3027 3022 3012 1 2 ND2 $T=863660 739320 1 180 $X=861800 $Y=738940
X1965 3034 3017 3041 1 2 ND2 $T=864900 729240 0 0 $X=864900 $Y=728860
X1966 3027 3035 3058 1 2 ND2 $T=864900 739320 0 0 $X=864900 $Y=738940
X1967 3053 2991 3017 1 2 ND2 $T=868000 729240 0 180 $X=866140 $Y=723820
X1968 3058 3056 3012 1 2 ND2 $T=868000 739320 0 0 $X=868000 $Y=738940
X1969 2935 3076 3044 1 2 ND2 $T=869860 880440 1 180 $X=868000 $Y=880060
X1970 3026 3064 3081 1 2 ND2 $T=870480 840120 1 0 $X=870480 $Y=834700
X1971 3066 3081 3054 1 2 ND2 $T=872960 840120 1 180 $X=871100 $Y=839740
X1972 3082 449 3072 1 2 ND2 $T=872960 729240 1 0 $X=872960 $Y=723820
X1973 3025 3103 3059 1 2 ND2 $T=875440 789720 1 180 $X=873580 $Y=789340
X1974 3088 3101 3071 1 2 ND2 $T=875440 860280 1 180 $X=873580 $Y=859900
X1975 3090 3108 3098 1 2 ND2 $T=877300 739320 1 180 $X=875440 $Y=738940
X1976 3118 3105 3075 1 2 ND2 $T=878540 779640 0 0 $X=878540 $Y=779260
X1977 3090 3119 3094 1 2 ND2 $T=879780 739320 0 0 $X=879780 $Y=738940
X1978 458 3124 456 1 2 ND2 $T=882880 900600 0 180 $X=881020 $Y=895180
X1979 3015 3161 3156 1 2 ND2 $T=884120 759480 0 0 $X=884120 $Y=759100
X1980 3115 3158 3163 1 2 ND2 $T=885360 789720 1 0 $X=885360 $Y=784300
X1981 3157 462 3180 1 2 ND2 $T=889080 729240 0 0 $X=889080 $Y=728860
X1982 3189 3183 3205 1 2 ND2 $T=891560 830040 1 0 $X=891560 $Y=824620
X1983 3222 3246 458 1 2 ND2 $T=897140 880440 1 0 $X=897140 $Y=875020
X1984 3208 3241 3240 1 2 ND2 $T=899000 739320 1 0 $X=899000 $Y=733900
X1985 3228 3251 3242 1 2 ND2 $T=903340 840120 0 180 $X=901480 $Y=834700
X1986 458 3274 3275 1 2 ND2 $T=905200 880440 1 0 $X=905200 $Y=875020
X1987 3331 3314 3301 1 2 ND2 $T=911400 799800 1 180 $X=909540 $Y=799420
X1988 3329 3308 3280 1 2 ND2 $T=913260 739320 0 0 $X=913260 $Y=738940
X1989 3147 490 494 1 2 ND2 $T=913880 900600 1 0 $X=913880 $Y=895180
X1990 3326 3356 3272 1 2 ND2 $T=914500 759480 1 0 $X=914500 $Y=754060
X1991 3371 3370 3376 1 2 ND2 $T=921940 830040 0 0 $X=921940 $Y=829660
X1992 3338 3371 3377 1 2 ND2 $T=921940 850200 1 0 $X=921940 $Y=844780
X1993 3415 3406 3400 1 2 ND2 $T=928140 850200 1 180 $X=926280 $Y=849820
X1994 3363 3411 3393 1 2 ND2 $T=928760 870360 1 180 $X=926900 $Y=869980
X1995 3272 3442 3422 1 2 ND2 $T=933720 759480 0 180 $X=931860 $Y=754060
X1996 3430 3444 3398 1 2 ND2 $T=933720 870360 0 180 $X=931860 $Y=864940
X1997 3438 3448 2798 1 2 ND2 $T=935580 799800 0 180 $X=933720 $Y=794380
X1998 3441 3467 3411 1 2 ND2 $T=936200 870360 1 180 $X=934340 $Y=869980
X1999 3444 3463 3411 1 2 ND2 $T=936820 870360 0 180 $X=934960 $Y=864940
X2000 3459 3478 3454 1 2 ND2 $T=936820 860280 1 0 $X=936820 $Y=854860
X2001 3439 3487 3459 1 2 ND2 $T=939920 850200 1 180 $X=938060 $Y=849820
X2002 3478 3481 3470 1 2 ND2 $T=942400 860280 0 180 $X=940540 $Y=854860
X2003 3456 3493 2744 1 2 ND2 $T=944880 779640 0 180 $X=943020 $Y=774220
X2004 3449 3510 3498 1 2 ND2 $T=946740 870360 1 180 $X=944880 $Y=869980
X2005 528 3523 3496 1 2 ND2 $T=948600 890520 1 180 $X=946740 $Y=890140
X2006 3494 3522 3523 1 2 ND2 $T=949220 860280 0 0 $X=949220 $Y=859900
X2007 3543 3551 3488 1 2 ND2 $T=954180 749400 0 0 $X=954180 $Y=749020
X2008 3526 3553 3540 1 2 ND2 $T=955420 880440 1 0 $X=955420 $Y=875020
X2009 3550 3546 539 1 2 ND2 $T=955420 890520 0 0 $X=955420 $Y=890140
X2010 3563 3566 3280 1 2 ND2 $T=958520 739320 1 180 $X=956660 $Y=738940
X2011 3526 3585 3569 1 2 ND2 $T=959140 880440 1 0 $X=959140 $Y=875020
X2012 3527 3594 3571 1 2 ND2 $T=964100 759480 1 180 $X=962240 $Y=759100
X2013 3526 3608 3575 1 2 ND2 $T=966580 870360 0 180 $X=964720 $Y=864940
X2014 3620 551 3632 1 2 ND2 $T=972780 729240 0 0 $X=972780 $Y=728860
X2015 3651 560 3652 1 2 ND2 $T=990760 749400 0 180 $X=988900 $Y=743980
X2016 695 687 1 669 2 664 OAI12HS $T=339760 769560 0 180 $X=336040 $Y=764140
X2017 679 626 1 676 2 697 OAI12HS $T=337280 799800 0 0 $X=337280 $Y=799420
X2018 720 722 1 707 2 687 OAI12HS $T=345340 759480 1 180 $X=341620 $Y=759100
X2019 721 742 1 715 2 698 OAI12HS $T=349060 729240 1 180 $X=345340 $Y=728860
X2020 730 734 1 736 2 735 OAI12HS $T=350920 799800 0 0 $X=350920 $Y=799420
X2021 732 693 1 703 2 716 OAI12HS $T=351540 749400 0 0 $X=351540 $Y=749020
X2022 763 753 1 728 2 715 OAI12HS $T=360220 729240 1 180 $X=356500 $Y=728860
X2023 778 786 1 791 2 714 OAI12HS $T=364560 809880 1 0 $X=364560 $Y=804460
X2024 817 795 1 777 2 791 OAI12HS $T=372000 799800 1 180 $X=368280 $Y=799420
X2025 38 849 1 856 2 794 OAI12HS $T=378820 729240 1 0 $X=378820 $Y=723820
X2026 1021 1015 1 1033 2 913 OAI12HS $T=417880 799800 0 0 $X=417880 $Y=799420
X2027 1056 1045 1 1002 2 1041 OAI12HS $T=423460 769560 0 180 $X=419740 $Y=764140
X2028 38 1088 1 1094 2 81 OAI12HS $T=431520 729240 1 0 $X=431520 $Y=723820
X2029 2422 332 1 2333 2 2446 OAI12HS $T=743380 749400 1 0 $X=743380 $Y=743980
X2030 2695 2590 1 2663 2 385 OAI12HS $T=801660 719160 0 0 $X=801660 $Y=718780
X2031 2789 2788 1 2805 2 2815 OAI12HS $T=821500 749400 1 0 $X=821500 $Y=743980
X2032 2784 403 1 2769 2 402 OAI12HS $T=827700 719160 1 180 $X=823980 $Y=718780
X2033 2769 2779 1 2803 2 2838 OAI12HS $T=824600 729240 1 0 $X=824600 $Y=723820
X2034 2871 2872 1 2885 2 2840 OAI12HS $T=836380 749400 1 0 $X=836380 $Y=743980
X2035 2870 414 1 2901 2 2915 OAI12HS $T=839480 890520 1 0 $X=839480 $Y=885100
X2036 3040 3048 1 3057 2 2992 OAI12HS $T=865520 779640 0 0 $X=865520 $Y=779260
X2037 3087 3048 1 3105 2 3099 OAI12HS $T=873580 769560 0 0 $X=873580 $Y=769180
X2038 414 3164 1 3124 2 3110 OAI12HS $T=884740 880440 0 180 $X=881020 $Y=875020
X2039 3149 3141 1 3078 2 3157 OAI12HS $T=887840 729240 1 180 $X=884120 $Y=728860
X2040 3185 3151 1 3159 2 3206 OAI12HS $T=895900 850200 0 180 $X=892180 $Y=844780
X2041 3238 3259 1 3241 2 479 OAI12HS $T=903340 729240 1 180 $X=899620 $Y=728860
X2042 478 3266 1 3246 2 3231 OAI12HS $T=903340 880440 0 180 $X=899620 $Y=875020
X2043 478 3264 1 3274 2 3273 OAI12HS $T=902720 870360 0 0 $X=902720 $Y=869980
X2044 3230 3162 1 3174 2 3299 OAI12HS $T=903340 789720 0 0 $X=903340 $Y=789340
X2045 3243 3193 1 3252 2 3281 OAI12HS $T=908300 860280 0 180 $X=904580 $Y=854860
X2046 3304 3295 1 485 2 3282 OAI12HS $T=910780 719160 1 180 $X=907060 $Y=718780
X2047 3300 3290 1 3281 2 3297 OAI12HS $T=911400 850200 0 180 $X=907680 $Y=844780
X2048 3257 3200 1 3308 2 3304 OAI12HS $T=908300 739320 0 0 $X=908300 $Y=738940
X2049 487 489 1 3282 2 497 OAI12HS $T=914500 719160 0 0 $X=914500 $Y=718780
X2050 3279 3382 1 3356 2 3357 OAI12HS $T=921320 759480 0 180 $X=917600 $Y=754060
X2051 3365 3334 1 3367 2 3368 OAI12HS $T=923800 860280 1 180 $X=920080 $Y=859900
X2052 3389 3403 1 3368 2 3400 OAI12HS $T=926280 860280 1 0 $X=926280 $Y=854860
X2053 3447 3279 1 3442 2 519 OAI12HS $T=938060 759480 0 180 $X=934340 $Y=754060
X2054 3547 3521 1 3566 2 3565 OAI12HS $T=957900 739320 1 0 $X=957900 $Y=733900
X2055 3555 3565 1 3518 2 3576 OAI12HS $T=965340 729240 1 180 $X=961620 $Y=728860
X2056 3586 3512 1 3594 2 3605 OAI12HS $T=964100 759480 1 0 $X=964100 $Y=754060
X2057 3598 3607 1 3576 2 3623 OAI12HS $T=967200 729240 0 0 $X=967200 $Y=728860
X2058 560 556 1 3638 2 558 OAI12HS $T=990140 719160 1 180 $X=986420 $Y=718780
X2059 610 627 1 634 2 NR2T $T=319920 749400 1 0 $X=319920 $Y=743980
X2060 638 596 1 624 2 NR2T $T=327360 769560 0 180 $X=322400 $Y=764140
X2061 18 698 1 694 2 NR2T $T=342240 729240 0 180 $X=337280 $Y=723820
X2062 3483 3449 1 3498 2 NR2T $T=939920 870360 0 0 $X=939920 $Y=869980
X2063 3499 528 1 3496 2 NR2T $T=949220 890520 0 180 $X=944260 $Y=885100
X2064 3554 3542 1 3487 2 NR2T $T=951700 850200 0 0 $X=951700 $Y=849820
X2065 3569 535 1 537 2 NR2T $T=954180 890520 1 0 $X=954180 $Y=885100
X2066 3575 3574 1 546 2 NR2T $T=964100 880440 0 0 $X=964100 $Y=880060
X2067 3622 546 1 3578 2 NR2T $T=967820 880440 1 0 $X=967820 $Y=875020
X2068 3625 3629 1 3622 2 NR2T $T=972780 880440 1 0 $X=972780 $Y=875020
X2069 559 3651 1 3652 2 NR2T $T=988280 739320 1 0 $X=988280 $Y=733900
X2070 612 1 11 597 2 616 ND3 $T=316820 739320 0 0 $X=316820 $Y=738940
X2071 628 1 625 606 2 618 ND3 $T=321780 789720 0 180 $X=319300 $Y=784300
X2072 638 1 623 621 2 11 ND3 $T=325500 799800 0 180 $X=323020 $Y=794380
X2073 640 1 638 618 2 11 ND3 $T=326740 789720 0 180 $X=324260 $Y=784300
X2074 646 1 649 655 2 662 ND3 $T=329220 779640 1 0 $X=329220 $Y=774220
X2075 638 1 647 667 2 11 ND3 $T=332320 789720 1 180 $X=329840 $Y=789340
X2076 638 1 631 662 2 13 ND3 $T=331080 769560 0 0 $X=331080 $Y=769180
X2077 2324 1 2441 2442 2 2330 ND3 $T=746480 759480 1 0 $X=746480 $Y=754060
X2078 2934 1 2925 2923 2 2917 ND3 $T=849400 870360 1 180 $X=846920 $Y=869980
X2079 3035 1 3022 3041 2 3056 ND3 $T=864900 739320 1 0 $X=864900 $Y=733900
X2080 3120 1 3119 3072 2 3108 ND3 $T=879780 739320 1 180 $X=877300 $Y=738940
X2081 3336 1 3171 3330 2 3293 ND3 $T=915740 830040 0 180 $X=913260 $Y=824620
X2082 3344 1 3330 3361 2 3325 ND3 $T=916360 819960 0 0 $X=916360 $Y=819580
X2083 3430 1 3467 3470 2 3475 ND3 $T=937440 870360 0 0 $X=937440 $Y=869980
X2084 3509 1 3541 3504 2 3428 ND3 $T=949840 840120 0 0 $X=949840 $Y=839740
X2085 3554 1 3540 3537 2 3414 ND3 $T=956040 870360 1 180 $X=953560 $Y=869980
X2086 3554 1 3569 3597 2 3414 ND3 $T=963480 870360 1 180 $X=961000 $Y=869980
X2087 3578 1 3585 3600 2 3597 ND3 $T=962860 880440 1 0 $X=962860 $Y=875020
X2088 590 593 7 2 1 XNR2HS $T=305040 739320 0 0 $X=305040 $Y=738940
X2089 651 644 14 2 1 XNR2HS $T=330460 729240 0 180 $X=324880 $Y=723820
X2090 669 665 629 2 1 XNR2HS $T=334180 769560 0 180 $X=328600 $Y=764140
X2091 13 657 15 2 1 XNR2HS $T=329840 719160 0 0 $X=329840 $Y=718780
X2092 663 678 656 2 1 XNR2HS $T=337280 749400 1 180 $X=331700 $Y=749020
X2093 703 701 666 2 1 XNR2HS $T=342860 749400 0 180 $X=337280 $Y=743980
X2094 682 688 678 2 1 XNR2HS $T=345340 759480 0 180 $X=339760 $Y=754060
X2095 695 687 665 2 1 XNR2HS $T=340380 769560 1 0 $X=340380 $Y=764140
X2096 720 725 663 2 1 XNR2HS $T=350920 759480 0 180 $X=345340 $Y=754060
X2097 734 729 708 2 1 XNR2HS $T=352780 789720 1 180 $X=347200 $Y=789340
X2098 738 737 684 2 1 XNR2HS $T=355260 779640 1 180 $X=349680 $Y=779260
X2099 730 736 729 2 1 XNR2HS $T=355880 799800 0 180 $X=350300 $Y=794380
X2100 744 740 732 2 1 XNR2HS $T=356500 759480 0 180 $X=350920 $Y=754060
X2101 748 743 724 2 1 XNR2HS $T=357120 749400 0 180 $X=351540 $Y=743980
X2102 764 761 703 2 1 XNR2HS $T=362080 759480 0 180 $X=356500 $Y=754060
X2103 768 760 743 2 1 XNR2HS $T=363320 749400 0 180 $X=357740 $Y=743980
X2104 739 745 737 2 1 XNR2HS $T=363320 779640 1 180 $X=357740 $Y=779260
X2105 777 773 705 2 1 XNR2HS $T=365180 799800 1 180 $X=359600 $Y=799420
X2106 769 783 682 2 1 XNR2HS $T=367040 759480 1 180 $X=361460 $Y=759100
X2107 772 797 763 2 1 XNR2HS $T=369520 749400 0 180 $X=363940 $Y=743980
X2108 788 787 22 2 1 XNR2HS $T=365800 729240 0 0 $X=365800 $Y=728860
X2109 803 822 736 2 1 XNR2HS $T=375720 799800 0 180 $X=370140 $Y=794380
X2110 782 789 761 2 1 XNR2HS $T=376960 759480 0 180 $X=371380 $Y=754060
X2111 795 817 773 2 1 XNR2HS $T=378200 799800 1 180 $X=372620 $Y=799420
X2112 833 828 806 2 1 XNR2HS $T=378820 769560 1 180 $X=373240 $Y=769180
X2113 834 775 798 2 1 XNR2HS $T=378820 779640 0 180 $X=373240 $Y=774220
X2114 845 830 801 2 1 XNR2HS $T=380680 749400 1 180 $X=375100 $Y=749020
X2115 832 805 822 2 1 XNR2HS $T=376340 799800 1 0 $X=376340 $Y=794380
X2116 826 810 36 2 1 XNR2HS $T=383160 739320 0 180 $X=377580 $Y=733900
X2117 868 866 719 2 1 XNR2HS $T=384400 799800 1 180 $X=378820 $Y=799420
X2118 878 829 843 2 1 XNR2HS $T=386260 789720 0 180 $X=380680 $Y=784300
X2119 902 899 795 2 1 XNR2HS $T=389980 799800 1 180 $X=384400 $Y=799420
X2120 851 46 862 2 1 XNR2HS $T=391840 749400 0 180 $X=386260 $Y=743980
X2121 878 841 855 2 1 XNR2HS $T=386880 789720 1 0 $X=386880 $Y=784300
X2122 830 892 41 2 1 XNR2HS $T=394320 739320 0 180 $X=388740 $Y=733900
X2123 830 912 49 2 1 XNR2HS $T=397420 729240 0 180 $X=391840 $Y=723820
X2124 940 929 718 2 1 XNR2HS $T=399280 779640 0 180 $X=393700 $Y=774220
X2125 946 851 930 2 1 XNR2HS $T=400520 769560 1 180 $X=394940 $Y=769180
X2126 920 913 899 2 1 XNR2HS $T=401140 799800 1 180 $X=395560 $Y=799420
X2127 912 965 925 2 1 XNR2HS $T=405480 749400 1 180 $X=399900 $Y=749020
X2128 975 974 959 2 1 XNR2HS $T=406720 789720 0 180 $X=401140 $Y=784300
X2129 965 53 934 2 1 XNR2HS $T=407340 749400 0 180 $X=401760 $Y=743980
X2130 959 977 868 2 1 XNR2HS $T=407340 799800 1 180 $X=401760 $Y=799420
X2131 56 973 911 2 1 XNR2HS $T=409200 739320 1 180 $X=403620 $Y=738940
X2132 981 833 994 2 1 XNR2HS $T=405480 789720 0 0 $X=405480 $Y=789340
X2133 1017 1001 939 2 1 XNR2HS $T=413540 729240 1 180 $X=407960 $Y=728860
X2134 976 827 1012 2 1 XNR2HS $T=410440 759480 0 0 $X=410440 $Y=759100
X2135 1017 1035 1007 2 1 XNR2HS $T=419740 739320 0 180 $X=414160 $Y=733900
X2136 981 841 1003 2 1 XNR2HS $T=420980 789720 0 180 $X=415400 $Y=784300
X2137 1002 1040 695 2 1 XNR2HS $T=421600 759480 1 180 $X=416020 $Y=759100
X2138 981 834 1013 2 1 XNR2HS $T=422840 789720 1 180 $X=417260 $Y=789340
X2139 70 1039 1015 2 1 XNR2HS $T=423460 769560 1 180 $X=417880 $Y=769180
X2140 981 829 1021 2 1 XNR2HS $T=423460 799800 0 180 $X=417880 $Y=794380
X2141 1045 1056 1040 2 1 XNR2HS $T=427800 759480 1 180 $X=422220 $Y=759100
X2142 1001 46 73 2 1 XNR2HS $T=424700 719160 0 0 $X=424700 $Y=718780
X2143 1073 968 1082 2 1 XNR2HS $T=427180 779640 1 0 $X=427180 $Y=774220
X2144 1001 84 86 2 1 XNR2HS $T=437100 729240 1 0 $X=437100 $Y=723820
X2145 1035 84 98 2 1 XNR2HS $T=448880 719160 0 0 $X=448880 $Y=718780
X2146 2199 279 280 2 1 XNR2HS $T=691300 729240 0 0 $X=691300 $Y=728860
X2147 291 2223 2257 2 1 XNR2HS $T=709280 729240 1 180 $X=703700 $Y=728860
X2148 291 2263 2271 2 1 XNR2HS $T=705560 739320 0 0 $X=705560 $Y=738940
X2149 2313 291 297 2 1 XNR2HS $T=717340 739320 1 180 $X=711760 $Y=738940
X2150 2324 2223 2336 2 1 XNR2HS $T=718580 769560 1 0 $X=718580 $Y=764140
X2151 2327 2223 2335 2 1 XNR2HS $T=726640 749400 0 180 $X=721060 $Y=743980
X2152 2327 2263 2374 2 1 XNR2HS $T=727880 739320 0 0 $X=727880 $Y=738940
X2153 290 2319 2377 2 1 XNR2HS $T=728500 749400 0 0 $X=728500 $Y=749020
X2154 2324 2263 2387 2 1 XNR2HS $T=731600 779640 1 0 $X=731600 $Y=774220
X2155 2355 320 333 2 1 XNR2HS $T=739040 729240 1 0 $X=739040 $Y=723820
X2156 299 2324 2422 2 1 XNR2HS $T=739660 759480 1 0 $X=739660 $Y=754060
X2157 2432 2424 2447 2 1 XNR2HS $T=744000 779640 1 0 $X=744000 $Y=774220
X2158 2256 2414 2451 2 1 XNR2HS $T=744620 739320 1 0 $X=744620 $Y=733900
X2159 2373 2451 2477 2 1 XNR2HS $T=750200 739320 1 0 $X=750200 $Y=733900
X2160 2458 2461 2478 2 1 XNR2HS $T=750200 769560 0 0 $X=750200 $Y=769180
X2161 2496 348 2520 2 1 XNR2HS $T=757640 729240 1 0 $X=757640 $Y=723820
X2162 2485 2478 2523 2 1 XNR2HS $T=758260 779640 1 0 $X=758260 $Y=774220
X2163 2434 2529 2551 2 1 XNR2HS $T=763220 759480 1 0 $X=763220 $Y=754060
X2164 2527 2568 2578 2 1 XNR2HS $T=767560 779640 1 0 $X=767560 $Y=774220
X2165 2401 2389 2586 2 1 XNR2HS $T=768800 759480 1 0 $X=768800 $Y=754060
X2166 2572 2580 2592 2 1 XNR2HS $T=770040 729240 0 0 $X=770040 $Y=728860
X2167 2551 2586 2610 2 1 XNR2HS $T=774380 759480 0 0 $X=774380 $Y=759100
X2168 2297 2538 2612 2 1 XNR2HS $T=775620 729240 0 0 $X=775620 $Y=728860
X2169 2283 2539 2613 2 1 XNR2HS $T=775620 739320 1 0 $X=775620 $Y=733900
X2170 2624 2585 2639 2 1 XNR2HS $T=789260 749400 1 180 $X=783680 $Y=749020
X2171 2641 2592 2679 2 1 XNR2HS $T=790500 729240 0 0 $X=790500 $Y=728860
X2172 2288 2562 2695 2 1 XNR2HS $T=794220 729240 1 0 $X=794220 $Y=723820
X2173 2704 2709 2731 2 1 XNR2HS $T=801660 759480 1 0 $X=801660 $Y=754060
X2174 2776 2768 2746 2 1 XNR2HS $T=820880 850200 0 180 $X=815300 $Y=844780
X2175 2810 400 2786 2 1 XNR2HS $T=825220 890520 0 180 $X=819640 $Y=885100
X2176 2801 2786 2809 2 1 XNR2HS $T=822120 880440 0 0 $X=822120 $Y=880060
X2177 2840 2844 406 2 1 XNR2HS $T=828940 739320 0 0 $X=828940 $Y=738940
X2178 2869 2876 2846 2 1 XNR2HS $T=838240 870360 0 180 $X=832660 $Y=864940
X2179 417 416 2870 2 1 XNR2HS $T=838860 890520 0 180 $X=833280 $Y=885100
X2180 2855 2882 419 2 1 XNR2HS $T=836380 729240 0 0 $X=836380 $Y=728860
X2181 2898 2896 2824 2 1 XNR2HS $T=842580 880440 0 180 $X=837000 $Y=875020
X2182 2907 421 2893 2 1 XNR2HS $T=844440 860280 1 180 $X=838860 $Y=859900
X2183 2890 2909 2833 2 1 XNR2HS $T=845680 850200 0 180 $X=840100 $Y=844780
X2184 2916 2913 2791 2 1 XNR2HS $T=846920 769560 0 180 $X=841340 $Y=764140
X2185 2911 2915 2898 2 1 XNR2HS $T=848160 880440 0 180 $X=842580 $Y=875020
X2186 2949 427 2801 2 1 XNR2HS $T=851880 890520 0 180 $X=846300 $Y=885100
X2187 2970 2967 2896 2 1 XNR2HS $T=855600 890520 1 180 $X=850020 $Y=890140
X2188 3010 436 2961 2 1 XNR2HS $T=863040 719160 1 180 $X=857460 $Y=718780
X2189 441 3037 2996 2 1 XNR2HS $T=866760 850200 1 180 $X=861180 $Y=849820
X2190 3006 2696 3040 2 1 XNR2HS $T=862420 789720 1 0 $X=862420 $Y=784300
X2191 3049 3019 3037 2 1 XNR2HS $T=870480 860280 0 180 $X=864900 $Y=854860
X2192 3071 3065 3049 2 1 XNR2HS $T=871100 860280 1 180 $X=865520 $Y=859900
X2193 398 443 3062 2 1 XNR2HS $T=865520 890520 0 0 $X=865520 $Y=890140
X2194 429 443 3089 2 1 XNR2HS $T=869860 890520 1 0 $X=869860 $Y=885100
X2195 3006 2683 3087 2 1 XNR2HS $T=877920 779640 1 180 $X=872340 $Y=779260
X2196 453 3110 3093 2 1 XNR2HS $T=878540 860280 0 180 $X=872960 $Y=854860
X2197 3101 3093 3100 2 1 XNR2HS $T=874200 850200 0 0 $X=874200 $Y=849820
X2198 3099 3074 3090 2 1 XNR2HS $T=874820 749400 1 0 $X=874820 $Y=743980
X2199 416 3111 3127 2 1 XNR2HS $T=876060 890520 1 0 $X=876060 $Y=885100
X2200 3078 3131 3113 2 1 XNR2HS $T=883500 729240 1 180 $X=877920 $Y=728860
X2201 3117 2683 3136 2 1 XNR2HS $T=877920 769560 1 0 $X=877920 $Y=764140
X2202 459 3126 3097 2 1 XNR2HS $T=884740 840120 1 180 $X=879160 $Y=839740
X2203 3149 3141 3131 2 1 XNR2HS $T=885360 739320 0 180 $X=879780 $Y=733900
X2204 3044 2935 3144 2 1 XNR2HS $T=879780 880440 0 0 $X=879780 $Y=880060
X2205 2744 3170 3153 2 1 XNR2HS $T=889700 769560 1 180 $X=884120 $Y=769180
X2206 463 3175 3159 2 1 XNR2HS $T=890320 850200 1 180 $X=884740 $Y=849820
X2207 437 3111 3178 2 1 XNR2HS $T=885360 890520 0 0 $X=885360 $Y=890140
X2208 3183 3171 3165 2 1 XNR2HS $T=891560 830040 0 180 $X=885980 $Y=824620
X2209 3159 3166 3181 2 1 XNR2HS $T=885980 840120 0 0 $X=885980 $Y=839740
X2210 3185 3151 3166 2 1 XNR2HS $T=892180 850200 0 180 $X=886600 $Y=844780
X2211 3148 3176 3185 2 1 XNR2HS $T=887220 860280 0 0 $X=887220 $Y=859900
X2212 3182 2741 3197 2 1 XNR2HS $T=889700 759480 1 0 $X=889700 $Y=754060
X2213 3187 3212 467 2 1 XNR2HS $T=896520 729240 0 180 $X=890940 $Y=723820
X2214 3182 2820 3186 2 1 XNR2HS $T=890940 759480 0 0 $X=890940 $Y=759100
X2215 2935 437 3209 2 1 XNR2HS $T=890940 880440 0 0 $X=890940 $Y=880060
X2216 438 3111 3202 2 1 XNR2HS $T=890940 900600 1 0 $X=890940 $Y=895180
X2217 3170 3198 3215 2 1 XNR2HS $T=892180 769560 0 0 $X=892180 $Y=769180
X2218 454 476 3247 2 1 XNR2HS $T=896520 900600 1 0 $X=896520 $Y=895180
X2219 475 3237 3252 2 1 XNR2HS $T=897140 860280 1 0 $X=897140 $Y=854860
X2220 3231 3218 3237 2 1 XNR2HS $T=897140 860280 0 0 $X=897140 $Y=859900
X2221 3258 3256 477 2 1 XNR2HS $T=903340 729240 0 180 $X=897760 $Y=723820
X2222 3236 3239 3253 2 1 XNR2HS $T=897760 819960 0 0 $X=897760 $Y=819580
X2223 454 480 3264 2 1 XNR2HS $T=899620 880440 0 0 $X=899620 $Y=880060
X2224 447 476 3270 2 1 XNR2HS $T=900240 890520 0 0 $X=900240 $Y=890140
X2225 3292 3287 484 2 1 XNR2HS $T=908920 729240 1 180 $X=903340 $Y=728860
X2226 3273 3262 3284 2 1 XNR2HS $T=903340 870360 1 0 $X=903340 $Y=864940
X2227 3276 2683 3289 2 1 XNR2HS $T=904580 779640 0 0 $X=904580 $Y=779260
X2228 2792 3276 3296 2 1 XNR2HS $T=905200 789720 1 0 $X=905200 $Y=784300
X2229 3255 3284 3324 2 1 XNR2HS $T=908920 860280 0 0 $X=908920 $Y=859900
X2230 3306 3225 3321 2 1 XNR2HS $T=909540 870360 0 0 $X=909540 $Y=869980
X2231 3294 3320 3319 2 1 XNR2HS $T=911400 850200 1 0 $X=911400 $Y=844780
X2232 3343 2798 3257 2 1 XNR2HS $T=917600 749400 1 180 $X=912020 $Y=749020
X2233 3332 3335 491 2 1 XNR2HS $T=918220 729240 0 180 $X=912640 $Y=723820
X2234 3357 3352 3335 2 1 XNR2HS $T=919460 739320 0 180 $X=913880 $Y=733900
X2235 3322 493 3359 2 1 XNR2HS $T=915120 870360 1 0 $X=915120 $Y=864940
X2236 3276 3198 3364 2 1 XNR2HS $T=916360 789720 1 0 $X=916360 $Y=784300
X2237 3365 3334 3351 2 1 XNR2HS $T=921940 860280 0 180 $X=916360 $Y=854860
X2238 3343 2813 3373 2 1 XNR2HS $T=917600 749400 0 0 $X=917600 $Y=749020
X2239 3367 3351 3377 2 1 XNR2HS $T=919460 850200 0 0 $X=919460 $Y=849820
X2240 2798 3353 3384 2 1 XNR2HS $T=920080 759480 0 0 $X=920080 $Y=759100
X2241 3370 3361 3385 2 1 XNR2HS $T=920080 819960 0 0 $X=920080 $Y=819580
X2242 3339 3359 3367 2 1 XNR2HS $T=920700 870360 1 0 $X=920700 $Y=864940
X2243 3393 3363 3378 2 1 XNR2HS $T=926280 870360 1 180 $X=920700 $Y=869980
X2244 3360 3381 505 2 1 XNR2HS $T=921320 729240 0 0 $X=921320 $Y=728860
X2245 3409 2741 3395 2 1 XNR2HS $T=929380 779640 0 180 $X=923800 $Y=774220
X2246 3316 2685 3405 2 1 XNR2HS $T=925660 759480 0 0 $X=925660 $Y=759100
X2247 3278 3345 3417 2 1 XNR2HS $T=925660 890520 0 0 $X=925660 $Y=890140
X2248 3398 3378 3415 2 1 XNR2HS $T=926280 870360 1 0 $X=926280 $Y=864940
X2249 3433 3397 512 2 1 XNR2HS $T=933720 729240 1 180 $X=928140 $Y=728860
X2250 3417 3431 3416 2 1 XNR2HS $T=933720 880440 0 180 $X=928140 $Y=875020
X2251 3409 2820 3423 2 1 XNR2HS $T=929380 779640 1 0 $X=929380 $Y=774220
X2252 515 3429 3440 2 1 XNR2HS $T=930620 860280 1 0 $X=930620 $Y=854860
X2253 3409 2685 3443 2 1 XNR2HS $T=931240 779640 0 0 $X=931240 $Y=779260
X2254 506 3418 3434 2 1 XNR2HS $T=931240 890520 0 0 $X=931240 $Y=890140
X2255 3316 2813 3447 2 1 XNR2HS $T=931860 759480 0 0 $X=931860 $Y=759100
X2256 3458 3455 518 2 1 XNR2HS $T=938060 719160 1 180 $X=932480 $Y=718780
X2257 3432 3414 3457 2 1 XNR2HS $T=933100 840120 1 0 $X=933100 $Y=834700
X2258 3434 3416 3464 2 1 XNR2HS $T=934340 880440 1 0 $X=934340 $Y=875020
X2259 3448 3462 3477 2 1 XNR2HS $T=936200 799800 1 0 $X=936200 $Y=794380
X2260 3465 3469 524 2 1 XNR2HS $T=937440 729240 0 0 $X=937440 $Y=728860
X2261 3445 3484 3472 2 1 XNR2HS $T=943640 799800 1 180 $X=938060 $Y=799420
X2262 3445 3340 3520 2 1 XNR2HS $T=944880 809880 1 0 $X=944880 $Y=804460
X2263 3456 2816 3524 2 1 XNR2HS $T=945500 779640 1 0 $X=945500 $Y=774220
X2264 3445 3503 3525 2 1 XNR2HS $T=945500 799800 0 0 $X=945500 $Y=799420
X2265 3488 3466 3530 2 1 XNR2HS $T=947360 749400 1 0 $X=947360 $Y=743980
X2266 3316 3466 3532 2 1 XNR2HS $T=947360 769560 1 0 $X=947360 $Y=764140
X2267 3445 3466 3533 2 1 XNR2HS $T=947360 789720 0 0 $X=947360 $Y=789340
X2268 3522 3506 3534 2 1 XNR2HS $T=947980 840120 1 0 $X=947980 $Y=834700
X2269 3340 3479 3536 2 1 XNR2HS $T=948600 769560 0 0 $X=948600 $Y=769180
X2270 3518 3548 3531 2 1 XNR2HS $T=956040 729240 1 180 $X=950460 $Y=728860
X2271 3488 3340 3547 2 1 XNR2HS $T=950460 739320 0 0 $X=950460 $Y=738940
X2272 3479 3503 3562 2 1 XNR2HS $T=954180 769560 0 0 $X=954180 $Y=769180
X2273 3555 3565 3548 2 1 XNR2HS $T=961620 729240 1 180 $X=956040 $Y=728860
X2274 3484 3479 3583 2 1 XNR2HS $T=959760 779640 1 0 $X=959760 $Y=774220
X2275 3477 3564 3590 2 1 XNR2HS $T=960380 799800 1 0 $X=960380 $Y=794380
X2276 3590 3573 548 2 1 XNR2HS $T=964720 789720 1 0 $X=964720 $Y=784300
X2277 3618 3600 3604 2 1 XNR2HS $T=972160 870360 1 180 $X=966580 $Y=869980
X2278 3626 3605 3615 2 1 XNR2HS $T=974020 759480 0 180 $X=968440 $Y=754060
X2279 3493 3451 3626 2 1 XNR2HS $T=977740 759480 1 180 $X=972160 $Y=759100
X2280 3630 3637 3643 2 1 XNR2HS $T=979600 769560 0 0 $X=979600 $Y=769180
X2281 3636 3634 3632 2 1 XNR2HS $T=980220 759480 1 0 $X=980220 $Y=754060
X2282 3616 3643 3651 2 1 XNR2HS $T=985180 769560 0 0 $X=985180 $Y=769180
X2283 3059 3025 3075 1 2 XOR2H $T=868000 789720 1 0 $X=868000 $Y=784300
X2284 3179 3196 3230 1 2 XOR2H $T=891560 799800 1 0 $X=891560 $Y=794380
X2285 624 2 613 596 1 NR2 $T=321160 769560 0 180 $X=319300 $Y=764140
X2286 639 2 611 633 1 NR2 $T=324880 799800 0 0 $X=324880 $Y=799420
X2287 666 2 635 674 1 NR2 $T=333560 739320 1 0 $X=333560 $Y=733900
X2288 672 2 683 628 1 NR2 $T=335420 799800 1 0 $X=335420 $Y=794380
X2289 697 2 685 683 1 NR2 $T=339760 799800 0 180 $X=337900 $Y=794380
X2290 706 2 679 714 1 NR2 $T=341620 809880 1 0 $X=341620 $Y=804460
X2291 739 2 746 738 1 NR2 $T=358980 789720 1 0 $X=358980 $Y=784300
X2292 769 2 759 774 1 NR2 $T=362080 769560 1 0 $X=362080 $Y=764140
X2293 747 2 758 731 1 NR2 $T=363320 739320 0 0 $X=363320 $Y=738940
X2294 772 2 748 779 1 NR2 $T=363320 749400 0 0 $X=363320 $Y=749020
X2295 810 2 776 819 1 NR2 $T=370760 739320 1 0 $X=370760 $Y=733900
X2296 805 2 813 803 1 NR2 $T=374480 789720 0 0 $X=374480 $Y=789340
X2297 38 2 869 875 1 NR2 $T=383160 729240 1 0 $X=383160 $Y=723820
X2298 855 2 888 850 1 NR2 $T=385640 799800 0 180 $X=383780 $Y=794380
X2299 837 2 907 915 1 NR2 $T=393700 789720 1 0 $X=393700 $Y=784300
X2300 986 2 926 978 1 NR2 $T=407960 779640 0 180 $X=406100 $Y=774220
X2301 978 2 987 985 1 NR2 $T=406100 779640 0 0 $X=406100 $Y=779260
X2302 62 2 979 978 1 NR2 $T=416640 779640 0 180 $X=414780 $Y=774220
X2303 58 2 1011 960 1 NR2 $T=415400 719160 0 0 $X=415400 $Y=718780
X2304 1035 2 1008 1025 1 NR2 $T=418500 739320 0 0 $X=418500 $Y=738940
X2305 1049 2 66 1015 1 NR2 $T=421600 749400 1 180 $X=419740 $Y=749020
X2306 1025 2 1045 1049 1 NR2 $T=419740 759480 1 0 $X=419740 $Y=754060
X2307 70 2 1065 1039 1 NR2 $T=425320 779640 1 0 $X=425320 $Y=774220
X2308 1072 2 1117 955 1 NR2 $T=440200 749400 1 180 $X=438340 $Y=749020
X2309 1035 2 1153 955 1 NR2 $T=449500 739320 0 180 $X=447640 $Y=733900
X2310 1153 2 1157 1114 1 NR2 $T=448260 729240 0 0 $X=448260 $Y=728860
X2311 1099 2 106 75 1 NR2 $T=461280 719160 0 0 $X=461280 $Y=718780
X2312 2195 2 2244 2235 1 NR2 $T=701220 729240 0 0 $X=701220 $Y=728860
X2313 2263 2 2242 2258 1 NR2 $T=705560 739320 1 0 $X=705560 $Y=733900
X2314 2282 2 2298 298 1 NR2 $T=711760 759480 1 0 $X=711760 $Y=754060
X2315 2305 2 2323 2312 1 NR2 $T=717960 749400 0 0 $X=717960 $Y=749020
X2316 2305 2 302 2258 1 NR2 $T=718580 729240 1 0 $X=718580 $Y=723820
X2317 2331 2 2339 2235 1 NR2 $T=721060 739320 1 0 $X=721060 $Y=733900
X2318 2334 2 310 2258 1 NR2 $T=725400 729240 1 0 $X=725400 $Y=723820
X2319 2258 2 330 2408 1 NR2 $T=739040 729240 0 0 $X=739040 $Y=728860
X2320 2408 2 2445 295 1 NR2 $T=744620 729240 0 0 $X=744620 $Y=728860
X2321 2441 2 2458 323 1 NR2 $T=748960 759480 1 0 $X=748960 $Y=754060
X2322 2263 2 2473 326 1 NR2 $T=750820 729240 0 0 $X=750820 $Y=728860
X2323 344 2 2493 326 1 NR2 $T=755780 729240 1 180 $X=753920 $Y=728860
X2324 2424 2 2502 2432 1 NR2 $T=755780 779640 0 180 $X=753920 $Y=774220
X2325 2441 2 2494 332 1 NR2 $T=757640 759480 1 180 $X=755780 $Y=759100
X2326 2482 2 2507 2495 1 NR2 $T=760120 779640 1 180 $X=758260 $Y=779260
X2327 2473 2 2522 2528 1 NR2 $T=761360 739320 1 0 $X=761360 $Y=733900
X2328 342 2 2531 2441 1 NR2 $T=762600 749400 1 0 $X=762600 $Y=743980
X2329 2494 2 2540 2511 1 NR2 $T=763220 769560 0 0 $X=763220 $Y=769180
X2330 2557 2 2568 2507 1 NR2 $T=766940 779640 0 0 $X=766940 $Y=779260
X2331 2445 2 2564 2446 1 NR2 $T=768180 739320 0 0 $X=768180 $Y=738940
X2332 2559 2 2588 2573 1 NR2 $T=769420 759480 0 0 $X=769420 $Y=759100
X2333 2539 2 2572 2581 1 NR2 $T=770040 739320 1 0 $X=770040 $Y=733900
X2334 2423 2 2603 2514 1 NR2 $T=776240 749400 1 0 $X=776240 $Y=743980
X2335 2538 2 361 2605 1 NR2 $T=778100 729240 1 0 $X=778100 $Y=723820
X2336 2599 2 2631 2627 1 NR2 $T=780580 779640 1 0 $X=780580 $Y=774220
X2337 2612 2 2638 2427 1 NR2 $T=781820 729240 1 0 $X=781820 $Y=723820
X2338 2640 2 2681 2662 1 NR2 $T=792980 759480 0 180 $X=791120 $Y=754060
X2339 2562 2 375 2675 1 NR2 $T=791740 719160 0 0 $X=791740 $Y=718780
X2340 2700 2 2713 2693 1 NR2 $T=800420 739320 1 180 $X=798560 $Y=738940
X2341 2692 2 2709 2681 1 NR2 $T=798560 759480 1 0 $X=798560 $Y=754060
X2342 2761 2 2756 2713 1 NR2 $T=817160 739320 0 0 $X=817160 $Y=738940
X2343 2764 2 2768 2767 1 NR2 $T=817160 840120 0 0 $X=817160 $Y=839740
X2344 2758 2 2779 2790 1 NR2 $T=819020 729240 0 0 $X=819020 $Y=728860
X2345 2780 2 2784 2797 1 NR2 $T=820260 739320 1 0 $X=820260 $Y=733900
X2346 2806 2 2788 2781 1 NR2 $T=823360 759480 0 180 $X=821500 $Y=754060
X2347 2779 2 2847 2784 1 NR2 $T=825840 729240 0 0 $X=825840 $Y=728860
X2348 400 2 2826 2810 1 NR2 $T=827080 890520 0 0 $X=827080 $Y=890140
X2349 2864 2 2868 2846 1 NR2 $T=835760 860280 1 180 $X=833900 $Y=859900
X2350 2866 2 2875 2868 1 NR2 $T=835140 860280 1 0 $X=835140 $Y=854860
X2351 2862 2 2837 413 1 NR2 $T=835140 880440 0 0 $X=835140 $Y=880060
X2352 2742 2 2872 2880 1 NR2 $T=835760 749400 0 0 $X=835760 $Y=749020
X2353 2900 2 2862 414 1 NR2 $T=840720 880440 1 180 $X=838860 $Y=880060
X2354 2904 2 2909 2879 1 NR2 $T=844440 850200 0 0 $X=844440 $Y=849820
X2355 426 2 2897 2900 1 NR2 $T=848160 870360 0 180 $X=846300 $Y=864940
X2356 2922 2 2889 2933 1 NR2 $T=847540 850200 0 0 $X=847540 $Y=849820
X2357 2927 2 2926 2942 1 NR2 $T=848780 759480 1 0 $X=848780 $Y=754060
X2358 2930 2 2913 2943 1 NR2 $T=848780 769560 0 0 $X=848780 $Y=769180
X2359 2931 2 2930 2944 1 NR2 $T=848780 779640 1 0 $X=848780 $Y=774220
X2360 2960 2 2969 2956 1 NR2 $T=853120 749400 1 0 $X=853120 $Y=743980
X2361 2977 2 2947 2969 1 NR2 $T=856220 739320 1 180 $X=854360 $Y=738940
X2362 2981 2 2984 2999 1 NR2 $T=856840 830040 0 0 $X=856840 $Y=829660
X2363 2998 2 2986 2987 1 NR2 $T=859320 769560 0 180 $X=857460 $Y=764140
X2364 433 2 2985 2972 1 NR2 $T=860560 860280 0 180 $X=858700 $Y=854860
X2365 3005 2 2952 3015 1 NR2 $T=860560 749400 0 0 $X=860560 $Y=749020
X2366 3002 2 3032 435 1 NR2 $T=863660 890520 1 180 $X=861800 $Y=890140
X2367 3014 2 2964 3000 1 NR2 $T=862420 759480 0 0 $X=862420 $Y=759100
X2368 3029 2 2937 2938 1 NR2 $T=864280 860280 1 180 $X=862420 $Y=859900
X2369 430 2 3002 3033 1 NR2 $T=862420 900600 1 0 $X=862420 $Y=895180
X2370 398 2 3029 442 1 NR2 $T=864900 880440 0 0 $X=864900 $Y=880060
X2371 3085 2 3078 3074 1 NR2 $T=872960 749400 0 180 $X=871100 $Y=743980
X2372 3015 2 3014 3083 1 NR2 $T=871720 759480 1 0 $X=871720 $Y=754060
X2373 3109 2 2974 3018 1 NR2 $T=877300 759480 0 180 $X=875440 $Y=754060
X2374 3009 2 3107 442 1 NR2 $T=877920 870360 1 180 $X=876060 $Y=869980
X2375 3059 2 3115 3025 1 NR2 $T=876680 789720 1 0 $X=876680 $Y=784300
X2376 453 2 3112 3110 1 NR2 $T=878540 860280 1 180 $X=876680 $Y=859900
X2377 3044 2 3104 2935 1 NR2 $T=877920 880440 0 0 $X=877920 $Y=880060
X2378 3116 2 3123 450 1 NR2 $T=877920 890520 0 0 $X=877920 $Y=890140
X2379 3138 2 3134 3123 1 NR2 $T=882260 890520 1 180 $X=880400 $Y=890140
X2380 3126 2 3130 459 1 NR2 $T=881020 850200 0 0 $X=881020 $Y=849820
X2381 3033 2 3138 3127 1 NR2 $T=884740 890520 1 180 $X=882880 $Y=890140
X2382 3140 2 3154 3134 1 NR2 $T=884740 860280 0 0 $X=884740 $Y=859900
X2383 3163 2 3173 3103 1 NR2 $T=889080 789720 0 180 $X=887220 $Y=784300
X2384 3089 2 3190 450 1 NR2 $T=888460 890520 1 0 $X=888460 $Y=885100
X2385 3196 2 3210 3170 1 NR2 $T=893420 789720 1 180 $X=891560 $Y=789340
X2386 3207 2 3224 3190 1 NR2 $T=895280 890520 0 180 $X=893420 $Y=885100
X2387 3202 2 3207 3033 1 NR2 $T=893420 890520 0 0 $X=893420 $Y=890140
X2388 3176 2 3218 3211 1 NR2 $T=895280 860280 0 0 $X=895280 $Y=859900
X2389 3198 2 3109 3086 1 NR2 $T=895900 759480 1 0 $X=895900 $Y=754060
X2390 3219 2 3255 3224 1 NR2 $T=897760 870360 0 0 $X=897760 $Y=869980
X2391 3069 2 3244 3086 1 NR2 $T=898380 749400 0 0 $X=898380 $Y=749020
X2392 3269 2 3236 3233 1 NR2 $T=903340 830040 0 180 $X=901480 $Y=824620
X2393 3172 2 3149 3271 1 NR2 $T=905820 759480 1 180 $X=903960 $Y=759100
X2394 3178 2 3285 470 1 NR2 $T=906440 890520 0 0 $X=906440 $Y=890140
X2395 3270 2 3310 486 1 NR2 $T=910780 890520 1 180 $X=908920 $Y=890140
X2396 3292 2 3332 3312 1 NR2 $T=912020 729240 0 0 $X=912020 $Y=728860
X2397 3310 2 3348 3285 1 NR2 $T=912020 890520 1 0 $X=912020 $Y=885100
X2398 3174 2 3337 3314 1 NR2 $T=914500 799800 0 180 $X=912640 $Y=794380
X2399 3306 2 3339 3315 1 NR2 $T=915120 880440 0 180 $X=913260 $Y=875020
X2400 3198 2 3333 3346 1 NR2 $T=914500 769560 1 0 $X=914500 $Y=764140
X2401 3321 2 3327 3294 1 NR2 $T=915740 860280 0 0 $X=915740 $Y=859900
X2402 3354 2 3358 3337 1 NR2 $T=918220 799800 0 180 $X=916360 $Y=794380
X2403 3325 2 3375 3347 1 NR2 $T=918840 840120 1 180 $X=916980 $Y=839740
X2404 3355 2 3369 3348 1 NR2 $T=918220 880440 0 0 $X=918220 $Y=880060
X2405 3346 2 3380 3172 1 NR2 $T=920700 769560 0 180 $X=918840 $Y=764140
X2406 3381 2 502 3362 1 NR2 $T=923800 729240 0 180 $X=921940 $Y=723820
X2407 3163 2 3396 3346 1 NR2 $T=925040 789720 1 0 $X=925040 $Y=784300
X2408 3345 2 507 3391 1 NR2 $T=927520 900600 0 180 $X=925660 $Y=895180
X2409 3249 2 3413 3346 1 NR2 $T=928760 779640 0 0 $X=928760 $Y=779260
X2410 3346 2 3427 3407 1 NR2 $T=931240 789720 0 180 $X=929380 $Y=784300
X2411 3400 2 3426 3415 1 NR2 $T=930000 850200 0 0 $X=930000 $Y=849820
X2412 3469 2 3508 3485 1 NR2 $T=943020 729240 1 0 $X=943020 $Y=723820
X2413 3417 2 3514 3431 1 NR2 $T=944880 880440 0 0 $X=944880 $Y=880060
X2414 526 2 3518 3500 1 NR2 $T=947980 729240 1 180 $X=946120 $Y=728860
X2415 3630 2 3645 3637 1 NR2 $T=982080 779640 0 0 $X=982080 $Y=779260
X2416 3644 2 556 3647 1 NR2 $T=983940 729240 1 0 $X=983940 $Y=723820
X2417 3640 2 3653 3639 1 NR2 $T=988900 769560 1 0 $X=988900 $Y=764140
X2418 636 2 642 1 627 NR2P $T=327360 739320 1 180 $X=323640 $Y=738940
X2419 632 2 629 1 603 NR2P $T=324880 759480 1 0 $X=324880 $Y=754060
X2420 641 2 637 1 599 NR2P $T=327360 759480 0 0 $X=327360 $Y=759100
X2421 650 2 633 1 623 NR2P $T=327360 799800 1 0 $X=327360 $Y=794380
X2422 650 2 672 1 647 NR2P $T=334800 799800 0 180 $X=331080 $Y=794380
X2423 652 2 656 1 636 NR2P $T=331700 749400 1 0 $X=331700 $Y=743980
X2424 712 2 708 1 691 NR2P $T=342240 789720 1 0 $X=342240 $Y=784300
X2425 709 2 705 1 633 NR2P $T=344100 799800 0 0 $X=344100 $Y=799420
X2426 787 2 790 1 731 NR2P $T=364560 739320 1 0 $X=364560 $Y=733900
X2427 2329 2 2258 1 303 NR2P $T=725400 729240 0 180 $X=721680 $Y=723820
X2428 314 2 2362 1 309 NR2P $T=729740 719160 1 180 $X=726020 $Y=718780
X2429 2355 2 2339 1 2362 NR2P $T=727880 729240 1 0 $X=727880 $Y=723820
X2430 314 2 2362 1 318 NR2P $T=734080 719160 1 180 $X=730360 $Y=718780
X2431 314 2 2362 1 329 NR2P $T=739040 719160 0 0 $X=739040 $Y=718780
X2432 2594 2 2579 1 2599 NR2P $T=772520 779640 0 0 $X=772520 $Y=779260
X2433 2804 2 2809 1 2762 NR2P $T=824600 870360 0 180 $X=820880 $Y=864940
X2434 2835 2 2839 1 2767 NR2P $T=827080 870360 1 0 $X=827080 $Y=864940
X2435 2899 2 2893 1 2879 NR2P $T=843820 860280 1 0 $X=843820 $Y=854860
X2436 2993 2 2982 1 2981 NR2P $T=856840 840120 0 0 $X=856840 $Y=839740
X2437 3139 2 3181 1 3199 NR2P $T=893420 840120 0 180 $X=889700 $Y=834700
X2438 3187 2 3227 1 471 NR2P $T=897760 719160 1 180 $X=894040 $Y=718780
X2439 3242 2 3228 1 3233 NR2P $T=897140 840120 1 0 $X=897140 $Y=834700
X2440 3232 2 3117 1 3204 NR2P $T=897760 789720 0 0 $X=897760 $Y=789340
X2441 3258 2 3286 1 485 NR2P $T=907680 729240 0 180 $X=903960 $Y=723820
X2442 3199 2 3233 1 3293 NR2P $T=907680 830040 0 0 $X=907680 $Y=829660
X2443 3297 2 3319 1 3311 NR2P $T=911400 840120 1 180 $X=907680 $Y=839740
X2444 3347 2 3311 1 3303 NR2P $T=915120 840120 1 0 $X=915120 $Y=834700
X2445 3338 2 3377 1 3347 NR2P $T=920700 850200 0 180 $X=916980 $Y=844780
X2446 3394 2 3375 1 3401 NR2P $T=925660 840120 1 180 $X=921940 $Y=839740
X2447 3433 2 3450 1 3455 NR2P $T=936820 729240 0 180 $X=933100 $Y=723820
X2448 3483 2 3499 1 3507 NR2P $T=947980 850200 1 180 $X=944260 $Y=849820
X2449 544 2 3606 1 3595 NR2P $T=966580 890520 1 180 $X=962860 $Y=890140
X2450 3578 2 3611 1 3606 NR2P $T=969060 890520 0 0 $X=969060 $Y=890140
X2451 738 739 1 746 712 751 2 MOAI1 $T=353400 789720 1 0 $X=353400 $Y=784300
X2452 775 26 1 785 752 793 2 MOAI1 $T=363320 789720 1 0 $X=363320 $Y=784300
X2453 26 784 1 785 762 800 2 MOAI1 $T=364560 779640 0 0 $X=364560 $Y=779260
X2454 26 812 1 785 765 798 2 MOAI1 $T=373240 769560 1 180 $X=368900 $Y=769180
X2455 803 805 1 813 777 821 2 MOAI1 $T=368900 789720 0 0 $X=368900 $Y=789340
X2456 26 815 1 801 747 31 2 MOAI1 $T=373860 739320 1 180 $X=369520 $Y=738940
X2457 26 825 1 31 34 41 2 MOAI1 $T=375100 719160 0 0 $X=375100 $Y=718780
X2458 840 37 1 850 749 860 2 MOAI1 $T=377580 759480 0 0 $X=377580 $Y=759100
X2459 864 854 1 843 754 837 2 MOAI1 $T=382540 779640 1 180 $X=378200 $Y=779260
X2460 863 37 1 850 782 853 2 MOAI1 $T=383780 759480 0 180 $X=379440 $Y=754060
X2461 44 921 1 910 48 38 2 MOAI1 $T=396180 719160 1 180 $X=391840 $Y=718780
X2462 942 941 1 937 783 930 2 MOAI1 $T=400520 769560 0 180 $X=396180 $Y=764140
X2463 942 998 1 937 766 1012 2 MOAI1 $T=409200 779640 1 0 $X=409200 $Y=774220
X2464 942 1008 1 917 60 1025 2 MOAI1 $T=409820 739320 0 0 $X=409820 $Y=738940
X2465 1052 1092 1 1099 80 1109 2 MOAI1 $T=432140 739320 1 0 $X=432140 $Y=733900
X2466 280 2242 1 287 2256 2258 2 MOAI1 $T=699980 739320 1 0 $X=699980 $Y=733900
X2467 2290 280 1 287 2283 2271 2 MOAI1 $T=714860 739320 0 180 $X=710520 $Y=733900
X2468 315 2368 1 2385 2401 2374 2 MOAI1 $T=732220 749400 1 0 $X=732220 $Y=743980
X2469 309 2347 1 2386 2395 323 2 MOAI1 $T=732840 729240 1 0 $X=732840 $Y=723820
X2470 309 322 1 323 324 327 2 MOAI1 $T=734080 719160 0 0 $X=734080 $Y=718780
X2471 2375 2330 1 2403 2434 2336 2 MOAI1 $T=735940 769560 1 0 $X=735940 $Y=764140
X2472 329 2368 1 323 2423 2335 2 MOAI1 $T=738420 749400 1 0 $X=738420 $Y=743980
X2473 2330 341 1 336 337 2450 2 MOAI1 $T=755160 719160 1 180 $X=750820 $Y=718780
X2474 2471 2393 1 342 2485 2490 2 MOAI1 $T=752060 759480 1 0 $X=752060 $Y=754060
X2475 2402 2471 1 342 2514 2521 2 MOAI1 $T=757640 749400 1 0 $X=757640 $Y=743980
X2476 2446 2445 1 2545 2550 2564 2 MOAI1 $T=763840 739320 0 0 $X=763840 $Y=738940
X2477 2612 2427 1 2638 368 2592 2 MOAI1 $T=786160 729240 1 0 $X=786160 $Y=723820
X2478 2810 400 1 2826 2814 2836 2 MOAI1 $T=825220 890520 1 0 $X=825220 $Y=885100
X2479 413 2862 1 2858 2804 2837 2 MOAI1 $T=834520 880440 0 180 $X=830180 $Y=875020
X2480 2953 2932 1 2979 2972 2990 2 MOAI1 $T=854360 860280 0 0 $X=854360 $Y=859900
X2481 3075 3061 1 3048 3012 3045 2 MOAI1 $T=871100 779640 0 180 $X=866760 $Y=774220
X2482 3132 3091 1 3005 3143 3150 2 MOAI1 $T=880400 749400 1 0 $X=880400 $Y=743980
X2483 3126 459 1 3100 3139 3130 2 MOAI1 $T=884740 850200 0 180 $X=880400 $Y=844780
X2484 3162 3156 1 3152 3094 3161 2 MOAI1 $T=890320 759480 1 180 $X=885980 $Y=759100
X2485 458 3167 1 414 3184 3209 2 MOAI1 $T=887840 880440 1 0 $X=887840 $Y=875020
X2486 451 483 1 470 3278 3247 2 MOAI1 $T=902720 900600 1 0 $X=902720 $Y=895180
X2487 3272 3288 1 3279 3295 3323 2 MOAI1 $T=907680 759480 1 0 $X=907680 $Y=754060
X2488 458 3291 1 478 3322 488 2 MOAI1 $T=907680 880440 0 0 $X=907680 $Y=880060
X2489 3294 3321 1 3327 3338 3324 2 MOAI1 $T=910780 860280 1 0 $X=910780 $Y=854860
X2490 3298 3333 1 3277 3208 3346 2 MOAI1 $T=913260 769560 0 0 $X=913260 $Y=769180
X2491 3298 3374 1 3277 3360 3296 2 MOAI1 $T=923180 769560 1 180 $X=918840 $Y=769180
X2492 3410 3408 1 3277 3397 3395 2 MOAI1 $T=930000 769560 1 180 $X=925660 $Y=769180
X2493 3452 3460 1 3451 3446 3005 2 MOAI1 $T=939300 749400 1 180 $X=934960 $Y=749020
X2494 3476 3410 1 3435 521 3443 2 MOAI1 $T=941160 779640 1 180 $X=936820 $Y=779260
X2495 3431 3417 1 3482 3498 3514 2 MOAI1 $T=941780 880440 1 0 $X=941780 $Y=875020
X2496 3527 3501 1 3512 3555 3532 2 MOAI1 $T=952940 769560 1 0 $X=952940 $Y=764140
X2497 3280 3570 1 3521 3591 3572 2 MOAI1 $T=961620 739320 0 0 $X=961620 $Y=738940
X2498 3527 3536 1 3602 3610 3512 2 MOAI1 $T=964720 759480 0 0 $X=964720 $Y=759100
X2499 3527 3562 1 3512 3628 3589 2 MOAI1 $T=966580 769560 0 0 $X=966580 $Y=769180
X2500 3630 3637 1 3645 3644 3648 2 MOAI1 $T=981460 779640 1 0 $X=981460 $Y=774220
X2501 640 1 620 625 2 ND2P $T=324260 779640 1 180 $X=320540 $Y=779260
X2502 631 1 620 649 2 ND2P $T=324880 779640 0 180 $X=321160 $Y=774220
X2503 623 1 620 619 2 ND2P $T=321160 789720 0 0 $X=321160 $Y=789340
X2504 647 1 620 670 2 ND2P $T=329840 789720 1 180 $X=326120 $Y=789340
X2505 666 1 674 642 2 ND2P $T=332940 739320 0 0 $X=332940 $Y=738940
X2506 2533 1 2610 2630 2 ND2P $T=780580 769560 0 180 $X=776860 $Y=764140
X2507 2630 1 2669 2656 2 ND2P $T=789260 769560 1 0 $X=789260 $Y=764140
X2508 2738 1 2713 2730 2 ND2P $T=809100 739320 1 0 $X=809100 $Y=733900
X2509 2796 1 2793 2823 2 ND2P $T=823980 840120 0 0 $X=823980 $Y=839740
X2510 2772 1 2766 2812 2 ND2P $T=823980 850200 0 0 $X=823980 $Y=849820
X2511 2804 1 2809 2772 2 ND2P $T=823980 860280 0 0 $X=823980 $Y=859900
X2512 2899 1 2893 2892 2 ND2P $T=843200 860280 0 180 $X=839480 $Y=854860
X2513 3017 1 2994 3020 2 ND2P $T=863040 729240 1 180 $X=859320 $Y=728860
X2514 2981 1 3026 3046 2 ND2P $T=869860 840120 1 180 $X=866140 $Y=839740
X2515 3139 1 3181 3205 2 ND2P $T=894040 830040 1 180 $X=890320 $Y=829660
X2516 3319 1 3297 3325 2 ND2P $T=915740 840120 1 180 $X=912020 $Y=839740
X2517 3261 1 3303 3392 2 ND2P $T=924420 840120 0 180 $X=920700 $Y=834700
X2518 3507 1 3481 3492 2 ND2P $T=947980 860280 0 180 $X=944260 $Y=854860
X2519 3577 1 3526 3582 2 ND2P $T=961620 860280 0 0 $X=961620 $Y=859900
X2520 3624 1 3613 547 2 ND2P $T=972160 719160 1 180 $X=968440 $Y=718780
X2521 704 711 718 1 2 677 MAO222 $T=346580 779640 0 180 $X=341620 $Y=774220
X2522 692 724 717 1 2 674 MAO222 $T=353400 739320 1 180 $X=348440 $Y=738940
X2523 760 748 768 1 2 693 MAO222 $T=362080 749400 1 180 $X=357120 $Y=749020
X2524 781 776 794 1 2 753 MAO222 $T=367040 729240 0 180 $X=362080 $Y=723820
X2525 782 764 789 1 2 688 MAO222 $T=367040 759480 0 180 $X=362080 $Y=754060
X2526 920 913 902 1 2 906 MAO222 $T=395560 799800 1 180 $X=390600 $Y=799420
X2527 901 929 955 1 2 739 MAO222 $T=400520 779640 1 180 $X=395560 $Y=779260
X2528 2256 2414 2373 1 2 2427 MAO222 $T=739660 739320 1 0 $X=739660 $Y=733900
X2529 2485 2461 2458 1 2 2533 MAO222 $T=753920 769560 1 0 $X=753920 $Y=764140
X2530 2395 2572 2469 1 2 2590 MAO222 $T=768800 729240 1 0 $X=768800 $Y=723820
X2531 2389 2551 2401 1 2 2633 MAO222 $T=775000 759480 1 0 $X=775000 $Y=754060
X2532 2550 2477 2613 1 2 2650 MAO222 $T=781820 739320 1 0 $X=781820 $Y=733900
X2533 3049 441 3019 1 2 3054 MAO222 $T=867380 850200 0 0 $X=867380 $Y=849820
X2534 463 3154 3184 1 2 3193 MAO222 $T=887220 860280 1 0 $X=887220 $Y=854860
X2535 3231 3218 475 1 2 3294 MAO222 $T=902720 860280 0 0 $X=902720 $Y=859900
X2536 3273 3255 482 1 2 3334 MAO222 $T=908920 870360 1 0 $X=908920 $Y=864940
X2537 3352 3332 3357 1 2 492 MAO222 $T=920080 729240 1 180 $X=915120 $Y=728860
X2538 3322 3339 493 1 2 3363 MAO222 $T=915120 870360 0 0 $X=915120 $Y=869980
X2539 3399 502 3387 1 2 513 MAO222 $T=925040 729240 1 0 $X=925040 $Y=723820
X2540 504 501 3369 1 2 3431 MAO222 $T=926900 880440 0 0 $X=926900 $Y=880060
X2541 3458 523 3455 1 2 530 MAO222 $T=939300 719160 0 0 $X=939300 $Y=718780
X2542 3601 3609 3612 1 2 3620 MAO222 $T=965960 739320 0 0 $X=965960 $Y=738940
X2543 3605 3493 3451 1 2 3609 MAO222 $T=974640 759480 1 0 $X=974640 $Y=754060
X2544 669 765 2 770 759 1 711 FA1 $T=350920 769560 0 0 $X=350920 $Y=769180
X2545 738 752 2 754 780 1 734 FA1 $T=368280 789720 1 180 $X=352780 $Y=789340
X2546 704 766 2 762 804 1 745 FA1 $T=371380 779640 0 180 $X=355880 $Y=774220
X2547 706 893 2 889 906 1 866 FA1 $T=376960 809880 1 0 $X=376960 $Y=804460
X2548 780 901 2 926 962 1 803 FA1 $T=404860 789720 1 180 $X=389360 $Y=789340
X2549 893 987 2 999 1022 1 977 FA1 $T=399900 809880 1 0 $X=399900 $Y=804460
X2550 3077 3145 2 3143 3113 1 465 FA1 $T=874820 719160 0 0 $X=874820 $Y=718780
X2551 3082 3145 2 3143 3113 1 3746 FA1 $T=874820 729240 1 0 $X=874820 $Y=723820
X2552 3449 529 2 525 520 1 3496 FA1 $T=935580 900600 1 0 $X=935580 $Y=895180
X2553 527 3544 2 3556 3508 1 3560 FA1 $T=946120 729240 1 0 $X=946120 $Y=723820
X2554 533 3560 2 3515 3531 1 540 FA1 $T=947360 719160 0 0 $X=947360 $Y=718780
X2555 3515 3446 2 3380 3519 1 3579 FA1 $T=947360 759480 1 0 $X=947360 $Y=754060
X2556 3647 3596 2 3299 3599 1 3573 FA1 $T=975880 789720 1 180 $X=960380 $Y=789340
X2557 542 3623 2 3615 3587 1 3624 FA1 $T=962860 729240 1 0 $X=962860 $Y=723820
X2558 3581 3493 2 3413 3545 1 3631 FA1 $T=962860 779640 0 0 $X=962860 $Y=779260
X2559 3587 3535 2 3591 3579 1 3612 FA1 $T=964720 749400 1 0 $X=964720 $Y=743980
X2560 3637 3557 2 3436 3621 1 3599 FA1 $T=981460 799800 0 180 $X=965960 $Y=794380
X2561 3639 3551 2 3628 3631 1 3616 FA1 $T=985180 769560 0 180 $X=969680 $Y=764140
X2562 3601 3614 2 3610 3581 1 3650 FA1 $T=972160 749400 0 0 $X=972160 $Y=749020
X2563 3640 3396 2 3633 3567 1 3630 FA1 $T=990760 789720 0 180 $X=975260 $Y=784300
X2564 633 679 2 1 672 OR2 $T=336660 799800 1 180 $X=334180 $Y=799420
X2565 688 682 2 1 671 OR2 $T=337900 759480 0 180 $X=335420 $Y=754060
X2566 755 740 2 1 720 OR2 $T=358980 759480 0 0 $X=358980 $Y=759100
X2567 888 907 2 1 902 OR2 $T=389980 799800 1 0 $X=389980 $Y=794380
X2568 991 1013 2 1 1033 OR2 $T=414780 799800 1 0 $X=414780 $Y=794380
X2569 1206 1157 2 1 111 OR2 $T=465000 719160 0 0 $X=465000 $Y=718780
X2570 2447 2454 2 1 2456 OR2 $T=751440 779640 1 180 $X=748960 $Y=779260
X2571 2536 2522 2 1 2560 OR2 $T=765080 769560 1 0 $X=765080 $Y=764140
X2572 2610 2533 2 1 2651 OR2 $T=782440 769560 1 0 $X=782440 $Y=764140
X2573 2639 2633 2 1 2647 OR2 $T=789260 759480 0 180 $X=786780 $Y=754060
X2574 2674 2664 2 1 2658 OR2 $T=792980 739320 1 180 $X=790500 $Y=738940
X2575 2824 2814 2 1 2787 OR2 $T=826460 870360 1 180 $X=823980 $Y=869980
X2576 2827 2817 2 1 2831 OR2 $T=831420 749400 1 180 $X=828940 $Y=749020
X2577 2830 2842 2 1 2853 OR2 $T=828940 860280 1 0 $X=828940 $Y=854860
X2578 421 2895 2 1 2864 OR2 $T=841960 870360 0 180 $X=839480 $Y=864940
X2579 2946 2937 2 1 2940 OR2 $T=851260 860280 1 0 $X=851260 $Y=854860
X2580 2968 2980 2 1 2957 OR2 $T=858080 779640 0 180 $X=855600 $Y=774220
X2581 2948 2986 2 1 2995 OR2 $T=856840 749400 1 0 $X=856840 $Y=743980
X2582 2978 2974 2 1 2936 OR2 $T=860560 759480 0 180 $X=858080 $Y=754060
X2583 3034 3041 2 1 3053 OR2 $T=870480 729240 1 180 $X=868000 $Y=728860
X2584 3077 3072 2 1 445 OR2 $T=871720 719160 1 180 $X=869240 $Y=718780
X2585 3214 3220 2 1 3240 OR2 $T=896520 739320 1 0 $X=896520 $Y=733900
X2586 486 3247 2 1 3328 OR2 $T=909540 900600 1 0 $X=909540 $Y=895180
X2587 3379 3342 2 1 506 OR2 $T=921940 890520 0 0 $X=921940 $Y=890140
X2588 3363 3393 2 1 3430 OR2 $T=928760 870360 0 0 $X=928760 $Y=869980
X2589 3463 3464 2 1 3459 OR2 $T=938060 870360 1 0 $X=938060 $Y=864940
X2590 3510 3499 2 1 3517 OR2 $T=946120 860280 0 0 $X=946120 $Y=859900
X2591 3629 546 2 1 3618 OR2 $T=973400 880440 1 180 $X=970920 $Y=880060
X2592 613 13 2 620 1 605 AOI12HS $T=317440 769560 0 0 $X=317440 $Y=769180
X2593 891 44 2 869 1 40 AOI12HS $T=387500 719160 1 180 $X=383160 $Y=718780
X2594 1001 1011 2 61 1 983 AOI12HS $T=410440 719160 0 0 $X=410440 $Y=718780
X2595 2223 2339 2 2355 1 2365 AOI12HS $T=726020 729240 0 0 $X=726020 $Y=728860
X2596 2735 2658 2 2713 1 2751 AOI12HS $T=811580 739320 0 0 $X=811580 $Y=738940
X2597 2840 2831 2 2818 1 2789 AOI12HS $T=830180 749400 0 180 $X=825840 $Y=743980
X2598 2815 2847 2 2838 1 409 AOI12HS $T=829560 729240 0 0 $X=829560 $Y=728860
X2599 2957 2916 2 2930 1 2929 AOI12HS $T=853120 769560 0 180 $X=848780 $Y=764140
X2600 3007 2823 2 2981 1 3028 AOI12HS $T=860560 830040 0 0 $X=860560 $Y=829660
X2601 2683 3204 2 3133 1 3226 AOI12HS $T=897760 779640 1 180 $X=893420 $Y=779260
X2602 3189 3171 2 3217 1 3239 AOI12HS $T=895900 830040 1 0 $X=895900 $Y=824620
X2603 3171 3293 2 3261 1 3302 AOI12HS $T=907060 830040 1 0 $X=907060 $Y=824620
X2604 3439 3428 2 3454 1 3461 AOI12HS $T=939920 850200 0 180 $X=935580 $Y=844780
X2605 3541 3428 2 3481 1 3491 AOI12HS $T=944880 840120 1 180 $X=940540 $Y=839740
X2606 3554 3414 2 3526 1 3561 AOI12HS $T=961000 860280 0 180 $X=956660 $Y=854860
X2607 609 605 9 2 1 XOR2HS $T=316820 769560 1 180 $X=311240 $Y=769180
X2608 601 608 12 2 1 XOR2HS $T=314340 729240 0 0 $X=314340 $Y=728860
X2609 704 702 641 2 1 XOR2HS $T=342860 769560 1 180 $X=337280 $Y=769180
X2610 710 693 701 2 1 XOR2HS $T=349680 749400 0 180 $X=344100 $Y=743980
X2611 718 711 702 2 1 XOR2HS $T=352780 779640 0 180 $X=347200 $Y=774220
X2612 749 733 725 2 1 XOR2HS $T=357740 759480 1 180 $X=352160 $Y=759100
X2613 829 775 812 2 1 XOR2HS $T=377580 779640 1 180 $X=372000 $Y=779260
X2614 830 827 815 2 1 XOR2HS $T=378200 749400 0 180 $X=372620 $Y=743980
X2615 831 828 816 2 1 XOR2HS $T=378200 769560 0 180 $X=372620 $Y=764140
X2616 841 775 784 2 1 XOR2HS $T=380060 789720 0 180 $X=374480 $Y=784300
X2617 851 830 825 2 1 XOR2HS $T=381300 739320 1 180 $X=375720 $Y=738940
X2618 878 892 844 2 1 XOR2HS $T=388740 739320 0 180 $X=383160 $Y=733900
X2619 827 878 863 2 1 XOR2HS $T=388740 759480 1 180 $X=383160 $Y=759100
X2620 878 834 854 2 1 XOR2HS $T=389980 779640 0 180 $X=384400 $Y=774220
X2621 831 46 846 2 1 XOR2HS $T=390600 769560 0 180 $X=385020 $Y=764140
X2622 845 46 853 2 1 XOR2HS $T=391840 749400 1 180 $X=386260 $Y=749020
X2623 912 46 875 2 1 XOR2HS $T=393700 729240 1 180 $X=388120 $Y=728860
X2624 833 915 857 2 1 XOR2HS $T=394940 769560 1 180 $X=389360 $Y=769180
X2625 960 53 891 2 1 XOR2HS $T=404240 719160 1 180 $X=398660 $Y=718780
X2626 968 901 940 2 1 XOR2HS $T=405480 779640 0 180 $X=399900 $Y=774220
X2627 960 973 921 2 1 XOR2HS $T=406720 729240 0 180 $X=401140 $Y=723820
X2628 965 892 950 2 1 XOR2HS $T=406720 759480 0 180 $X=401140 $Y=754060
X2629 976 845 941 2 1 XOR2HS $T=410440 759480 1 180 $X=404860 $Y=759100
X2630 981 831 998 2 1 XOR2HS $T=409820 769560 0 0 $X=409820 $Y=769180
X2631 1017 982 980 2 1 XOR2HS $T=419740 729240 0 180 $X=414160 $Y=723820
X2632 1039 982 72 2 1 XOR2HS $T=422840 729240 1 0 $X=422840 $Y=723820
X2633 1071 845 1059 2 1 XOR2HS $T=428420 749400 1 180 $X=422840 $Y=749020
X2634 1071 851 1044 2 1 XOR2HS $T=428420 759480 0 180 $X=422840 $Y=754060
X2635 1071 827 1079 2 1 XOR2HS $T=434000 749400 1 180 $X=428420 $Y=749020
X2636 968 833 1078 2 1 XOR2HS $T=434000 769560 1 180 $X=428420 $Y=769180
X2637 1039 1035 1098 2 1 XOR2HS $T=430900 729240 0 0 $X=430900 $Y=728860
X2638 968 829 1076 2 1 XOR2HS $T=437720 779640 1 180 $X=432140 $Y=779260
X2639 968 841 1086 2 1 XOR2HS $T=438340 779640 0 180 $X=432760 $Y=774220
X2640 968 831 1083 2 1 XOR2HS $T=440200 769560 1 180 $X=434620 $Y=769180
X2641 1132 912 1092 2 1 XOR2HS $T=442680 739320 0 180 $X=437100 $Y=733900
X2642 1132 892 1050 2 1 XOR2HS $T=442680 739320 1 180 $X=437100 $Y=738940
X2643 84 973 85 2 1 XOR2HS $T=443300 719160 1 180 $X=437720 $Y=718780
X2644 1132 53 1125 2 1 XOR2HS $T=446400 729240 1 180 $X=440820 $Y=728860
X2645 84 982 1146 2 1 XOR2HS $T=443300 729240 1 0 $X=443300 $Y=723820
X2646 973 90 1183 2 1 XOR2HS $T=454460 719160 0 0 $X=454460 $Y=718780
X2647 90 1001 1191 2 1 XOR2HS $T=454460 729240 0 0 $X=454460 $Y=728860
X2648 1132 982 1224 2 1 XOR2HS $T=464380 729240 0 0 $X=464380 $Y=728860
X2649 291 2276 2290 2 1 XOR2HS $T=708660 749400 1 0 $X=708660 $Y=743980
X2650 298 2282 2330 2 1 XOR2HS $T=716720 759480 0 0 $X=716720 $Y=759100
X2651 2235 2313 2347 2 1 XOR2HS $T=721060 739320 0 0 $X=721060 $Y=738940
X2652 2319 289 312 2 1 XOR2HS $T=722920 739320 1 0 $X=722920 $Y=733900
X2653 2223 298 2360 2 1 XOR2HS $T=724780 759480 0 0 $X=724780 $Y=759100
X2654 2327 2276 2368 2 1 XOR2HS $T=726640 749400 1 0 $X=726640 $Y=743980
X2655 2324 2313 2375 2 1 XOR2HS $T=727880 769560 1 0 $X=727880 $Y=764140
X2656 2313 2382 2393 2 1 XOR2HS $T=732220 759480 0 0 $X=732220 $Y=759100
X2657 290 2382 2402 2 1 XOR2HS $T=734080 749400 0 0 $X=734080 $Y=749020
X2658 2276 2324 2407 2 1 XOR2HS $T=735320 769560 0 0 $X=735320 $Y=769180
X2659 2276 2382 2416 2 1 XOR2HS $T=738420 759480 0 0 $X=738420 $Y=759100
X2660 288 2382 2439 2 1 XOR2HS $T=742760 739320 0 0 $X=742760 $Y=738940
X2661 2355 288 2450 2 1 XOR2HS $T=744620 729240 1 0 $X=744620 $Y=723820
X2662 299 2382 2467 2 1 XOR2HS $T=748340 749400 0 0 $X=748340 $Y=749020
X2663 296 2382 2470 2 1 XOR2HS $T=748960 739320 0 0 $X=748960 $Y=738940
X2664 2445 2446 2571 2 1 XOR2HS $T=766320 749400 1 0 $X=766320 $Y=743980
X2665 2545 2571 2585 2 1 XOR2HS $T=768800 749400 0 0 $X=768800 $Y=749020
X2666 2395 2469 2580 2 1 XOR2HS $T=770660 719160 0 0 $X=770660 $Y=718780
X2667 2560 2587 2597 2 1 XOR2HS $T=771280 769560 1 0 $X=771280 $Y=764140
X2668 2514 2423 2624 2 1 XOR2HS $T=778100 749400 0 0 $X=778100 $Y=749020
X2669 2612 2427 2641 2 1 XOR2HS $T=781820 729240 0 0 $X=781820 $Y=728860
X2670 2613 2550 2646 2 1 XOR2HS $T=782440 739320 0 0 $X=782440 $Y=738940
X2671 2547 2631 2670 2 1 XOR2HS $T=787400 779640 1 0 $X=787400 $Y=774220
X2672 2477 2646 2674 2 1 XOR2HS $T=788640 739320 1 0 $X=788640 $Y=733900
X2673 2669 2710 2723 2 1 XOR2HS $T=799800 769560 1 0 $X=799800 $Y=764140
X2674 2695 2590 2727 2 1 XOR2HS $T=801040 729240 1 0 $X=801040 $Y=723820
X2675 2663 2727 391 2 1 XOR2HS $T=807240 719160 0 0 $X=807240 $Y=718780
X2676 2750 2751 394 2 1 XOR2HS $T=812820 729240 1 0 $X=812820 $Y=723820
X2677 2735 2756 2763 2 1 XOR2HS $T=813440 739320 1 0 $X=813440 $Y=733900
X2678 2766 2794 2774 2 1 XOR2HS $T=823980 850200 1 180 $X=818400 $Y=849820
X2679 2789 2808 404 2 1 XOR2HS $T=822740 739320 0 0 $X=822740 $Y=738940
X2680 2863 2875 2852 2 1 XOR2HS $T=838240 850200 0 180 $X=832660 $Y=844780
X2681 417 398 411 2 1 XOR2HS $T=838860 900600 0 180 $X=833280 $Y=895180
X2682 2862 413 2876 2 1 XOR2HS $T=835140 870360 0 0 $X=835140 $Y=869980
X2683 2936 2928 2905 2 1 XOR2HS $T=850640 759480 1 180 $X=845060 $Y=759100
X2684 2929 2947 2924 2 1 XOR2HS $T=852500 739320 1 180 $X=846920 $Y=738940
X2685 2940 2965 2903 2 1 XOR2HS $T=855600 850200 0 180 $X=850020 $Y=844780
X2686 2951 416 2953 2 1 XOR2HS $T=851260 880440 0 0 $X=851260 $Y=880060
X2687 2951 429 2941 2 1 XOR2HS $T=851880 880440 1 0 $X=851880 $Y=875020
X2688 2992 2987 2968 2 1 XOR2HS $T=859320 769560 1 180 $X=853740 $Y=769180
X2689 2994 2991 2962 2 1 XOR2HS $T=859940 729240 0 180 $X=854360 $Y=723820
X2690 3002 435 2970 2 1 XOR2HS $T=861180 900600 0 180 $X=855600 $Y=895180
X2691 438 434 2988 2 1 XOR2HS $T=863040 880440 1 180 $X=857460 $Y=880060
X2692 2823 2984 2989 2 1 XOR2HS $T=864280 830040 0 180 $X=858700 $Y=824620
X2693 3027 3023 2948 2 1 XOR2HS $T=865520 749400 0 180 $X=859940 $Y=743980
X2694 3025 2744 3008 2 1 XOR2HS $T=865520 769560 1 180 $X=859940 $Y=769180
X2695 3006 2744 3021 2 1 XOR2HS $T=859940 779640 1 0 $X=859940 $Y=774220
X2696 434 437 2997 2 1 XOR2HS $T=859940 880440 1 0 $X=859940 $Y=875020
X2697 3064 3028 2971 2 1 XOR2HS $T=870480 830040 0 180 $X=864900 $Y=824620
X2698 3058 3012 3023 2 1 XOR2HS $T=871100 749400 0 180 $X=865520 $Y=743980
X2699 3025 2792 3039 2 1 XOR2HS $T=871100 769560 1 180 $X=865520 $Y=769180
X2700 444 443 3067 2 1 XOR2HS $T=866140 900600 1 0 $X=866140 $Y=895180
X2701 3051 447 3060 2 1 XOR2HS $T=872960 880440 0 180 $X=867380 $Y=875020
X2702 3094 3090 3073 2 1 XOR2HS $T=875440 739320 1 180 $X=869860 $Y=738940
X2703 3098 3073 3034 2 1 XOR2HS $T=876060 739320 0 180 $X=870480 $Y=733900
X2704 2683 3095 3047 2 1 XOR2HS $T=876060 769560 0 180 $X=870480 $Y=764140
X2705 3100 3097 3066 2 1 XOR2HS $T=876060 850200 0 180 $X=870480 $Y=844780
X2706 3095 2820 3068 2 1 XOR2HS $T=877920 759480 1 180 $X=872340 $Y=759100
X2707 3051 454 3092 2 1 XOR2HS $T=881020 880440 0 180 $X=875440 $Y=875020
X2708 3095 2741 3091 2 1 XOR2HS $T=883500 759480 0 180 $X=877920 $Y=754060
X2709 3134 3140 3126 2 1 XOR2HS $T=884120 860280 1 180 $X=878540 $Y=859900
X2710 3095 2798 3169 2 1 XOR2HS $T=884120 759480 1 0 $X=884120 $Y=754060
X2711 3179 2792 3118 2 1 XOR2HS $T=890320 779640 1 180 $X=884740 $Y=779260
X2712 3051 464 3160 2 1 XOR2HS $T=890320 870360 1 180 $X=884740 $Y=869980
X2713 438 2935 3167 2 1 XOR2HS $T=885360 880440 0 0 $X=885360 $Y=880060
X2714 3194 3208 466 2 1 XOR2HS $T=895900 739320 0 180 $X=890320 $Y=733900
X2715 3154 3192 3175 2 1 XOR2HS $T=890940 850200 0 0 $X=890940 $Y=849820
X2716 3051 468 3203 2 1 XOR2HS $T=890940 870360 0 0 $X=890940 $Y=869980
X2717 3220 3214 3194 2 1 XOR2HS $T=897140 739320 1 180 $X=891560 $Y=738940
X2718 3224 3219 3243 2 1 XOR2HS $T=896520 870360 1 0 $X=896520 $Y=864940
X2719 3252 3254 3228 2 1 XOR2HS $T=903340 850200 0 180 $X=897760 $Y=844780
X2720 3193 3243 3254 2 1 XOR2HS $T=897760 850200 0 0 $X=897760 $Y=849820
X2721 3117 2792 3234 2 1 XOR2HS $T=904580 769560 1 180 $X=899000 $Y=769180
X2722 2685 3229 3191 2 1 XOR2HS $T=907060 749400 0 180 $X=901480 $Y=743980
X2723 480 447 3275 2 1 XOR2HS $T=905200 890520 1 0 $X=905200 $Y=885100
X2724 3305 3302 3263 2 1 XOR2HS $T=911400 819960 1 180 $X=905820 $Y=819580
X2725 3229 2813 3283 2 1 XOR2HS $T=912020 749400 1 180 $X=906440 $Y=749020
X2726 2816 3229 3313 2 1 XOR2HS $T=907680 749400 1 0 $X=907680 $Y=743980
X2727 3316 2820 3288 2 1 XOR2HS $T=913260 759480 1 180 $X=907680 $Y=759100
X2728 3276 2744 3317 2 1 XOR2HS $T=916360 789720 0 180 $X=910780 $Y=784300
X2729 3321 3324 3320 2 1 XOR2HS $T=916360 850200 1 180 $X=910780 $Y=849820
X2730 2741 3353 3323 2 1 XOR2HS $T=919460 759480 1 180 $X=913880 $Y=759100
X2731 3343 2685 3329 2 1 XOR2HS $T=920080 749400 0 180 $X=914500 $Y=743980
X2732 3348 3355 3365 2 1 XOR2HS $T=916360 880440 1 0 $X=916360 $Y=875020
X2733 3387 3386 500 2 1 XOR2HS $T=925660 719160 1 180 $X=920080 $Y=718780
X2734 2821 3265 3372 2 1 XOR2HS $T=926280 749400 0 180 $X=920700 $Y=743980
X2735 3369 501 3390 2 1 XOR2HS $T=920700 880440 0 0 $X=920700 $Y=880060
X2736 3342 3379 3393 2 1 XOR2HS $T=920700 890520 1 0 $X=920700 $Y=885100
X2737 504 3390 3398 2 1 XOR2HS $T=922560 880440 1 0 $X=922560 $Y=875020
X2738 3170 3383 3404 2 1 XOR2HS $T=923800 799800 0 0 $X=923800 $Y=799420
X2739 3343 2816 3412 2 1 XOR2HS $T=926280 749400 0 0 $X=926280 $Y=749020
X2740 3343 2821 3421 2 1 XOR2HS $T=926900 749400 1 0 $X=926900 $Y=743980
X2741 517 516 3418 2 1 XOR2HS $T=933720 900600 0 180 $X=928140 $Y=895180
X2742 3466 3265 3424 2 1 XOR2HS $T=939300 749400 0 180 $X=933720 $Y=743980
X2743 2798 3445 3408 2 1 XOR2HS $T=933720 789720 0 0 $X=933720 $Y=789340
X2744 3474 3461 3453 2 1 XOR2HS $T=940540 840120 1 180 $X=934960 $Y=839740
X2745 3340 3265 3437 2 1 XOR2HS $T=942400 739320 1 180 $X=936820 $Y=738940
X2746 3456 2813 3476 2 1 XOR2HS $T=936820 789720 1 0 $X=936820 $Y=784300
X2747 3316 2816 3480 2 1 XOR2HS $T=937440 759480 0 0 $X=937440 $Y=759100
X2748 3503 3265 3486 2 1 XOR2HS $T=946740 749400 0 180 $X=941160 $Y=743980
X2749 3316 2821 3501 2 1 XOR2HS $T=941780 769560 1 0 $X=941780 $Y=764140
X2750 3490 3491 3502 2 1 XOR2HS $T=941780 840120 1 0 $X=941780 $Y=834700
X2751 3484 3265 3460 2 1 XOR2HS $T=949220 749400 1 180 $X=943640 $Y=749020
X2752 2821 3456 3516 2 1 XOR2HS $T=944260 779640 0 0 $X=944260 $Y=779260
X2753 3488 3503 3563 2 1 XOR2HS $T=954800 749400 1 0 $X=954800 $Y=743980
X2754 3558 3561 3568 2 1 XOR2HS $T=956040 850200 1 0 $X=956040 $Y=844780
X2755 3488 3484 3570 2 1 XOR2HS $T=956660 749400 0 0 $X=956660 $Y=749020
X2756 3484 3479 3589 2 1 XOR2HS $T=960380 769560 0 0 $X=960380 $Y=769180
X2757 552 3627 3619 2 1 XOR2HS $T=974640 860280 1 180 $X=969060 $Y=859900
X2758 3640 3639 3634 2 1 XOR2HS $T=983320 759480 1 180 $X=977740 $Y=759100
X2759 816 26 1 31 811 760 2 MOAI1S $T=373860 749400 1 180 $X=370140 $Y=749020
X2760 864 862 1 853 852 768 2 MOAI1S $T=383160 749400 0 180 $X=379440 $Y=743980
X2761 864 908 1 837 903 929 2 MOAI1S $T=390600 779640 0 0 $X=390600 $Y=779260
X2762 37 921 1 983 989 57 2 MOAI1S $T=405480 719160 0 0 $X=405480 $Y=718780
X2763 981 942 1 991 1003 974 2 MOAI1S $T=407960 789720 1 0 $X=407960 $Y=784300
X2764 1183 1114 1 1099 1148 95 2 MOAI1S $T=453220 729240 0 180 $X=449500 $Y=723820
X2765 99 1191 1 1101 1209 109 2 MOAI1S $T=460040 729240 0 0 $X=460040 $Y=728860
X2766 2347 315 1 2338 2365 2373 2 MOAI1S $T=734700 729240 1 180 $X=730980 $Y=728860
X2767 2360 2465 1 2505 2509 2511 2 MOAI1S $T=756400 759480 1 0 $X=756400 $Y=754060
X2768 2514 2423 1 2585 2603 2664 2 MOAI1S $T=779340 749400 1 0 $X=779340 $Y=743980
X2769 2976 2941 1 426 2963 2869 2 MOAI1S $T=856220 870360 1 180 $X=852500 $Y=869980
X2770 3018 3039 1 3005 3036 3027 2 MOAI1S $T=868000 749400 1 180 $X=864280 $Y=749020
X2771 2976 2997 1 426 3050 2911 2 MOAI1S $T=864280 870360 0 0 $X=864280 $Y=869980
X2772 3047 2920 1 3052 3030 3000 2 MOAI1S $T=869860 759480 1 180 $X=866140 $Y=759100
X2773 451 3067 1 450 3062 3071 2 MOAI1S $T=876060 900600 0 180 $X=872340 $Y=895180
X2774 3162 3153 1 3152 3136 3146 2 MOAI1S $T=887220 769560 0 180 $X=883500 $Y=764140
X2775 3158 3179 1 3173 3179 3177 2 MOAI1S $T=889080 789720 1 0 $X=889080 $Y=784300
X2776 3215 3162 1 3188 3152 3098 2 MOAI1S $T=895900 769560 0 180 $X=892180 $Y=764140
X2777 3162 3234 1 3152 3248 3245 2 MOAI1S $T=897760 759480 0 0 $X=897760 $Y=759100
X2778 3230 3234 1 3226 3235 3214 2 MOAI1S $T=901480 779640 0 180 $X=897760 $Y=774220
X2779 3412 3280 1 3200 3373 3387 2 MOAI1S $T=927520 739320 1 180 $X=923800 $Y=738940
X2780 3272 3384 1 3279 3405 3399 2 MOAI1S $T=925040 759480 1 0 $X=925040 $Y=754060
X2781 3280 3421 1 3200 3419 514 2 MOAI1S $T=934960 739320 1 180 $X=931240 $Y=738940
X2782 3272 3473 1 3279 3489 3458 2 MOAI1S $T=939920 759480 1 0 $X=939920 $Y=754060
X2783 3445 3410 1 3341 3472 3462 2 MOAI1S $T=946120 799800 0 180 $X=942400 $Y=794380
X2784 3410 3516 1 3435 3524 3535 2 MOAI1S $T=956660 779640 0 180 $X=952940 $Y=774220
X2785 3410 3539 1 3341 3520 3557 2 MOAI1S $T=953560 799800 1 0 $X=953560 $Y=794380
X2786 3410 3552 1 3341 3533 3567 2 MOAI1S $T=954180 789720 0 0 $X=954180 $Y=789340
X2787 3488 3280 1 3521 3588 3614 2 MOAI1S $T=962240 749400 0 0 $X=962240 $Y=749020
X2788 3527 3583 1 3479 3512 3621 2 MOAI1S $T=965960 779640 1 0 $X=965960 $Y=774220
X2789 642 657 661 2 1 ND2S $T=330460 729240 0 0 $X=330460 $Y=728860
X2790 681 643 675 2 1 ND2S $T=333560 779640 0 0 $X=333560 $Y=779260
X2791 723 709 735 2 1 ND2S $T=348440 799800 0 0 $X=348440 $Y=799420
X2792 785 820 30 2 1 ND2S $T=372000 759480 0 0 $X=372000 $Y=759100
X2793 88 89 1146 2 1 ND2S $T=443920 719160 0 0 $X=443920 $Y=718780
X2794 2511 2526 2494 2 1 ND2S $T=761980 769560 1 180 $X=760120 $Y=769180
X2795 2651 2710 2630 2 1 ND2S $T=799800 759480 1 180 $X=797940 $Y=759100
X2796 2738 2750 2712 2 1 ND2S $T=811580 729240 1 180 $X=809720 $Y=728860
X2797 2782 396 2769 2 1 ND2S $T=820880 719160 1 180 $X=819020 $Y=718780
X2798 2775 399 2803 2 1 ND2S $T=822120 729240 1 0 $X=822120 $Y=723820
X2799 2795 2808 2805 2 1 ND2S $T=823980 749400 0 0 $X=823980 $Y=749020
X2800 2900 2891 417 2 1 ND2S $T=841960 890520 1 180 $X=840100 $Y=890140
X2801 2915 2934 2911 2 1 ND2S $T=850640 870360 0 0 $X=850640 $Y=869980
X2802 2950 2928 2959 2 1 ND2S $T=851260 759480 0 0 $X=851260 $Y=759100
X2803 2983 2965 2958 2 1 ND2S $T=857460 850200 1 180 $X=855600 $Y=849820
X2804 3000 2950 3014 2 1 ND2S $T=859320 759480 0 0 $X=859320 $Y=759100
X2805 3075 3057 3021 2 1 ND2S $T=871720 779640 1 180 $X=869860 $Y=779260
X2806 3094 3120 3098 2 1 ND2S $T=885360 739320 1 0 $X=885360 $Y=733900
X2807 3141 3180 3149 2 1 ND2S $T=887220 739320 1 0 $X=887220 $Y=733900
X2808 3325 3305 3336 2 1 ND2S $T=912640 819960 0 0 $X=912640 $Y=819580
X2809 3336 3344 3261 2 1 ND2S $T=916980 830040 1 0 $X=916980 $Y=824620
X2810 3438 3436 2820 2 1 ND2S $T=932480 799800 0 180 $X=930620 $Y=794380
X2811 3406 3432 3439 2 1 ND2S $T=931860 850200 1 0 $X=931860 $Y=844780
X2812 3459 3474 3470 2 1 ND2S $T=940540 860280 1 180 $X=938680 $Y=859900
X2813 3509 3490 3510 2 1 ND2S $T=946120 840120 0 0 $X=946120 $Y=839740
X2814 3521 3543 3195 2 1 ND2S $T=952320 749400 1 180 $X=950460 $Y=749020
X2815 3540 3558 534 2 1 ND2S $T=957280 870360 0 0 $X=957280 $Y=869980
X2816 3644 3638 3647 2 1 ND2S $T=987040 729240 1 180 $X=985180 $Y=728860
X2817 731 747 1 758 717 767 2 MOAI1H $T=354640 739320 0 0 $X=354640 $Y=738940
X2818 942 980 1 945 59 1007 2 MOAI1H $T=404860 739320 1 0 $X=404860 $Y=733900
X2819 407 410 1 414 2810 2891 2 MOAI1H $T=832660 890520 0 0 $X=832660 $Y=890140
X2820 3002 435 1 2967 3019 3032 2 MOAI1H $T=860560 890520 1 0 $X=860560 $Y=885100
X2821 3076 448 1 3104 450 448 2 MOAI1H $T=870480 880440 0 0 $X=870480 $Y=880060
X2822 453 3110 1 3101 3151 3112 2 MOAI1H $T=878540 860280 1 0 $X=878540 $Y=854860
X2823 3309 3298 1 3277 3256 3268 2 MOAI1H $T=910780 779640 0 180 $X=903340 $Y=774220
X2824 3298 3317 1 3341 3212 3364 2 MOAI1H $T=912020 779640 0 0 $X=912020 $Y=779260
X2825 3527 3480 1 3512 3556 3559 2 MOAI1H $T=951080 759480 0 0 $X=951080 $Y=759100
X2826 3639 3640 1 3653 3652 3636 2 MOAI1H $T=985800 759480 1 0 $X=985800 $Y=754060
X2827 13 622 1 2 INV2 $T=320540 729240 0 0 $X=320540 $Y=728860
X2828 650 640 1 2 INV2 $T=330460 789720 0 180 $X=328600 $Y=784300
X2829 691 675 1 2 INV2 $T=339760 789720 0 180 $X=337900 $Y=784300
X2830 753 742 1 2 INV2 $T=358360 729240 1 0 $X=358360 $Y=723820
X2831 797 779 1 2 INV2 $T=368280 749400 1 180 $X=366420 $Y=749020
X2832 788 790 1 2 INV2 $T=370140 739320 0 180 $X=368280 $Y=733900
X2833 37 873 1 2 INV2 $T=383160 749400 1 180 $X=381300 $Y=749020
X2834 864 850 1 2 INV2 $T=383160 779640 0 180 $X=381300 $Y=774220
X2835 870 38 1 2 INV2 $T=384400 729240 1 180 $X=382540 $Y=728860
X2836 873 870 1 2 INV2 $T=383780 749400 0 0 $X=383780 $Y=749020
X2837 870 837 1 2 INV2 $T=386880 769560 0 0 $X=386880 $Y=769180
X2838 897 44 1 2 INV2 $T=389360 719160 1 180 $X=387500 $Y=718780
X2839 897 864 1 2 INV2 $T=388120 729240 1 0 $X=388120 $Y=723820
X2840 933 942 1 2 INV2 $T=400520 769560 1 0 $X=400520 $Y=764140
X2841 967 933 1 2 INV2 $T=404860 769560 0 180 $X=403000 $Y=764140
X2842 954 923 1 2 INV2 $T=406100 890520 0 0 $X=406100 $Y=890140
X2843 996 917 1 2 INV2 $T=409820 749400 1 180 $X=407960 $Y=749020
X2844 961 981 1 2 INV2 $T=407960 769560 0 0 $X=407960 $Y=769180
X2845 996 945 1 2 INV2 $T=410440 749400 0 180 $X=408580 $Y=743980
X2846 954 1032 1 2 INV2 $T=415400 890520 0 0 $X=415400 $Y=890140
X2847 1015 967 1 2 INV2 $T=417880 769560 1 180 $X=416020 $Y=769180
X2848 1039 915 1 2 INV2 $T=419740 779640 0 180 $X=417880 $Y=774220
X2849 1034 897 1 2 INV2 $T=419740 729240 1 0 $X=419740 $Y=723820
X2850 1101 1052 1 2 INV2 $T=434620 749400 0 180 $X=432760 $Y=743980
X2851 1101 1075 1 2 INV2 $T=435240 759480 0 180 $X=433380 $Y=754060
X2852 1117 1101 1 2 INV2 $T=437100 749400 1 180 $X=435240 $Y=749020
X2853 1119 1131 1 2 INV2 $T=438340 779640 1 0 $X=438340 $Y=774220
X2854 1127 968 1 2 INV2 $T=440820 769560 0 180 $X=438960 $Y=764140
X2855 1132 955 1 2 INV2 $T=443920 749400 1 0 $X=443920 $Y=743980
X2856 1070 1119 1 2 INV2 $T=445780 789720 0 0 $X=445780 $Y=789340
X2857 1101 1114 1 2 INV2 $T=446400 739320 0 0 $X=446400 $Y=738940
X2858 1119 1154 1 2 INV2 $T=447640 789720 1 0 $X=447640 $Y=784300
X2859 1126 1213 1 2 INV2 $T=461900 850200 0 0 $X=461900 $Y=849820
X2860 1213 1226 1 2 INV2 $T=466240 860280 0 0 $X=466240 $Y=859900
X2861 132 1250 1 2 INV2 $T=492900 840120 0 0 $X=492900 $Y=839740
X2862 1369 127 1 2 INV2 $T=496620 739320 0 180 $X=494760 $Y=733900
X2863 1358 1282 1 2 INV2 $T=497860 799800 1 0 $X=497860 $Y=794380
X2864 1374 134 1 2 INV2 $T=500960 739320 1 180 $X=499100 $Y=738940
X2865 1443 1381 1 2 INV2 $T=515220 890520 0 180 $X=513360 $Y=885100
X2866 1459 1443 1 2 INV2 $T=520180 890520 0 180 $X=518320 $Y=885100
X2867 1447 1460 1 2 INV2 $T=522040 840120 1 0 $X=522040 $Y=834700
X2868 1460 1422 1 2 INV2 $T=522040 850200 1 0 $X=522040 $Y=844780
X2869 1504 1457 1 2 INV2 $T=528860 739320 1 180 $X=527000 $Y=738940
X2870 135 1468 1 2 INV2 $T=527000 749400 0 0 $X=527000 $Y=749020
X2871 132 1552 1 2 INV2 $T=540020 850200 0 0 $X=540020 $Y=849820
X2872 1646 1551 1 2 INV2 $T=556140 759480 1 180 $X=554280 $Y=759100
X2873 1561 1646 1 2 INV2 $T=562340 749400 0 0 $X=562340 $Y=749020
X2874 199 1796 1 2 INV2 $T=598920 870360 0 180 $X=597060 $Y=864940
X2875 1837 1840 1 2 INV2 $T=605740 759480 0 0 $X=605740 $Y=759100
X2876 135 1956 1 2 INV2 $T=616280 729240 0 0 $X=616280 $Y=728860
X2877 210 1504 1 2 INV2 $T=618140 739320 0 180 $X=616280 $Y=733900
X2878 234 1951 1 2 INV2 $T=638600 870360 1 0 $X=638600 $Y=864940
X2879 280 295 1 2 INV2 $T=713000 719160 0 0 $X=713000 $Y=718780
X2880 298 326 1 2 INV2 $T=736560 729240 0 0 $X=736560 $Y=728860
X2881 305 2403 1 2 INV2 $T=736560 759480 1 0 $X=736560 $Y=754060
X2882 2417 2280 1 2 INV2 $T=739660 819960 0 180 $X=737800 $Y=814540
X2883 305 336 1 2 INV2 $T=747100 719160 0 0 $X=747100 $Y=718780
X2884 2330 332 1 2 INV2 $T=754540 749400 1 0 $X=754540 $Y=743980
X2885 2493 2489 1 2 INV2 $T=755780 729240 0 0 $X=755780 $Y=728860
X2886 2489 2471 1 2 INV2 $T=756400 739320 0 0 $X=756400 $Y=738940
X2887 2489 352 1 2 INV2 $T=762600 719160 1 180 $X=760740 $Y=718780
X2888 2516 342 1 2 INV2 $T=761360 729240 0 0 $X=761360 $Y=728860
X2889 2523 2579 1 2 INV2 $T=772520 779640 1 180 $X=770660 $Y=779260
X2890 2635 2673 1 2 INV2 $T=791740 819960 1 0 $X=791740 $Y=814540
X2891 2681 2678 1 2 INV2 $T=795460 749400 1 180 $X=793600 $Y=749020
X2892 2628 2720 1 2 INV2 $T=799180 789720 0 0 $X=799180 $Y=789340
X2893 2706 2648 1 2 INV2 $T=799180 900600 1 0 $X=799180 $Y=895180
X2894 2720 2729 1 2 INV2 $T=802900 789720 0 0 $X=802900 $Y=789340
X2895 2720 2747 1 2 INV2 $T=807240 789720 0 0 $X=807240 $Y=789340
X2896 2767 2796 1 2 INV2 $T=821500 840120 0 0 $X=821500 $Y=839740
X2897 2762 2799 1 2 INV2 $T=825220 860280 1 0 $X=825220 $Y=854860
X2898 2417 2851 1 2 INV2 $T=827080 819960 1 0 $X=827080 $Y=814540
X2899 2886 2884 1 2 INV2 $T=838240 830040 0 180 $X=836380 $Y=824620
X2900 2886 2914 1 2 INV2 $T=843820 830040 1 0 $X=843820 $Y=824620
X2901 2906 2918 1 2 INV2 $T=846920 850200 1 0 $X=846920 $Y=844780
X2902 2996 2982 1 2 INV2 $T=858080 850200 0 180 $X=856220 $Y=844780
X2903 439 2899 1 2 INV2 $T=863660 860280 0 180 $X=861800 $Y=854860
X2904 2918 3051 1 2 INV2 $T=865520 880440 1 0 $X=865520 $Y=875020
X2905 3111 448 1 2 INV2 $T=876680 890520 1 180 $X=874820 $Y=890140
X2906 3121 3018 1 2 INV2 $T=879780 749400 1 180 $X=877920 $Y=749020
X2907 3107 3042 1 2 INV2 $T=879160 870360 0 0 $X=879160 $Y=869980
X2908 3042 3147 1 2 INV2 $T=881020 870360 0 0 $X=881020 $Y=869980
X2909 3033 451 1 2 INV2 $T=883500 900600 1 0 $X=883500 $Y=895180
X2910 3144 461 1 2 INV2 $T=885980 900600 1 0 $X=885980 $Y=895180
X2911 461 3033 1 2 INV2 $T=888460 900600 1 0 $X=888460 $Y=895180
X2912 3001 3133 1 2 INV2 $T=890320 779640 1 0 $X=890320 $Y=774220
X2913 3216 3250 1 2 INV2 $T=899000 789720 1 0 $X=899000 $Y=784300
X2914 3244 3121 1 2 INV2 $T=900240 749400 0 0 $X=900240 $Y=749020
X2915 3230 3152 1 2 INV2 $T=900240 769560 1 0 $X=900240 $Y=764140
X2916 3086 3265 1 2 INV2 $T=902100 749400 0 0 $X=902100 $Y=749020
X2917 3121 3267 1 2 INV2 $T=903340 739320 1 0 $X=903340 $Y=733900
X2918 3174 3350 1 2 INV2 $T=913880 789720 0 0 $X=913880 $Y=789340
X2919 3271 3298 1 2 INV2 $T=917600 779640 1 0 $X=917600 $Y=774220
X2920 3366 3341 1 2 INV2 $T=920700 789720 1 180 $X=918840 $Y=789340
X2921 3358 3366 1 2 INV2 $T=918840 799800 1 0 $X=918840 $Y=794380
X2922 3388 3276 1 2 INV2 $T=924420 789720 0 180 $X=922560 $Y=784300
X2923 3331 3388 1 2 INV2 $T=922560 799800 1 0 $X=922560 $Y=794380
X2924 3404 3402 1 2 INV2 $T=928140 799800 0 180 $X=926280 $Y=794380
X2925 3402 3271 1 2 INV2 $T=930000 789720 1 180 $X=928140 $Y=789340
X2926 3271 3410 1 2 INV2 $T=939920 789720 0 0 $X=939920 $Y=789340
X2927 3507 3542 1 2 INV2 $T=951700 860280 1 0 $X=951700 $Y=854860
X2928 549 3678 1 2 INV2 $T=1010600 719160 0 0 $X=1010600 $Y=718780
X2929 3681 3663 1 2 INV2 $T=1016180 749400 1 180 $X=1014320 $Y=749020
X2930 3680 3681 1 2 INV2 $T=1019280 749400 1 180 $X=1017420 $Y=749020
X2931 31 785 1 2 BUF2 $T=370760 759480 0 180 $X=367660 $Y=754060
X2932 824 886 1 2 BUF2 $T=393080 860280 1 0 $X=393080 $Y=854860
X2933 992 1090 1 2 BUF2 $T=430900 840120 0 0 $X=430900 $Y=839740
X2934 1110 1048 1 2 BUF2 $T=438960 819960 1 180 $X=435860 $Y=819580
X2935 1062 1072 1 2 BUF2 $T=437720 749400 1 0 $X=437720 $Y=743980
X2936 1090 1029 1 2 BUF2 $T=440820 830040 0 180 $X=437720 $Y=824620
X2937 1029 1070 1 2 BUF2 $T=438340 809880 1 0 $X=438340 $Y=804460
X2938 1048 1126 1 2 BUF2 $T=438960 840120 0 0 $X=438960 $Y=839740
X2939 90 1132 1 2 BUF2 $T=446400 739320 0 180 $X=443300 $Y=733900
X2940 99 1062 1 2 BUF2 $T=453840 729240 1 180 $X=450740 $Y=728860
X2941 1241 1172 1 2 BUF2 $T=473680 779640 1 180 $X=470580 $Y=779260
X2942 1238 1275 1 2 BUF2 $T=475540 830040 0 0 $X=475540 $Y=829660
X2943 100 1234 1 2 BUF2 $T=475540 890520 0 0 $X=475540 $Y=890140
X2944 1220 122 1 2 BUF2 $T=485460 729240 0 0 $X=485460 $Y=728860
X2945 1275 1293 1 2 BUF2 $T=494760 809880 1 0 $X=494760 $Y=804460
X2946 122 140 1 2 BUF2 $T=498480 719160 0 0 $X=498480 $Y=718780
X2947 1395 1447 1 2 BUF2 $T=519560 830040 0 0 $X=519560 $Y=829660
X2948 172 1459 1 2 BUF2 $T=545600 880440 1 180 $X=542500 $Y=880060
X2949 177 1382 1 2 BUF2 $T=551180 739320 0 180 $X=548080 $Y=733900
X2950 1622 172 1 2 BUF2 $T=560480 870360 1 180 $X=557380 $Y=869980
X2951 1653 1374 1 2 BUF2 $T=565440 739320 0 180 $X=562340 $Y=733900
X2952 1579 1669 1 2 BUF2 $T=565440 769560 0 0 $X=565440 $Y=769180
X2953 1635 1722 1 2 BUF2 $T=575980 759480 0 0 $X=575980 $Y=759100
X2954 1745 1647 1 2 BUF2 $T=586520 729240 1 180 $X=583420 $Y=728860
X2955 1358 199 1 2 BUF2 $T=593340 769560 1 0 $X=593340 $Y=764140
X2956 185 1751 1 2 BUF2 $T=593340 880440 0 0 $X=593340 $Y=880060
X2957 194 1826 1 2 BUF2 $T=603260 900600 1 0 $X=603260 $Y=895180
X2958 1798 1863 1 2 BUF2 $T=610080 759480 0 0 $X=610080 $Y=759100
X2959 1826 219 1 2 BUF2 $T=623720 900600 1 0 $X=623720 $Y=895180
X2960 1951 1982 1 2 BUF2 $T=639220 850200 0 0 $X=639220 $Y=849820
X2961 1982 1907 1 2 BUF2 $T=644800 830040 1 180 $X=641700 $Y=829660
X2962 1907 2012 1 2 BUF2 $T=647900 809880 0 180 $X=644800 $Y=804460
X2963 1956 2096 1 2 BUF2 $T=663400 739320 1 0 $X=663400 $Y=733900
X2964 2092 2078 1 2 BUF2 $T=675180 870360 1 180 $X=672080 $Y=869980
X2965 2096 275 1 2 BUF2 $T=685720 729240 1 0 $X=685720 $Y=723820
X2966 2227 2129 1 2 BUF2 $T=698120 840120 1 180 $X=695020 $Y=839740
X2967 279 2235 1 2 BUF2 $T=696880 739320 1 0 $X=696880 $Y=733900
X2968 2147 2219 1 2 BUF2 $T=696880 759480 0 0 $X=696880 $Y=759100
X2969 2147 2243 1 2 BUF2 $T=699360 769560 0 0 $X=699360 $Y=769180
X2970 2234 1589 1 2 BUF2 $T=699360 799800 0 0 $X=699360 $Y=799420
X2971 2265 2234 1 2 BUF2 $T=706180 809880 1 0 $X=706180 $Y=804460
X2972 2209 2267 1 2 BUF2 $T=713620 809880 1 180 $X=710520 $Y=809500
X2973 2267 2227 1 2 BUF2 $T=714860 840120 0 180 $X=711760 $Y=834700
X2974 2267 2320 1 2 BUF2 $T=714860 840120 1 0 $X=714860 $Y=834700
X2975 282 2265 1 2 BUF2 $T=718580 850200 0 0 $X=718580 $Y=849820
X2976 2319 2324 1 2 BUF2 $T=729740 759480 1 0 $X=729740 $Y=754060
X2977 2320 2378 1 2 BUF2 $T=729740 830040 1 0 $X=729740 $Y=824620
X2978 2433 2479 1 2 BUF2 $T=750200 789720 0 0 $X=750200 $Y=789340
X2979 2508 2435 1 2 BUF2 $T=769420 870360 0 180 $X=766320 $Y=864940
X2980 2589 2508 1 2 BUF2 $T=773760 880440 1 180 $X=770660 $Y=880060
X2981 2479 2628 1 2 BUF2 $T=780580 789720 1 0 $X=780580 $Y=784300
X2982 2619 2417 1 2 BUF2 $T=781200 819960 1 0 $X=781200 $Y=814540
X2983 2569 2660 1 2 BUF2 $T=788020 809880 0 0 $X=788020 $Y=809500
X2984 2661 376 1 2 BUF2 $T=802280 799800 1 0 $X=802280 $Y=794380
X2985 3174 3117 1 2 BUF2 $T=888460 789720 0 0 $X=888460 $Y=789340
X2986 3048 3200 1 2 BUF2 $T=895900 749400 0 180 $X=892800 $Y=743980
X2987 478 414 1 2 BUF2 $T=899620 880440 1 180 $X=896520 $Y=880060
X2988 3250 3272 1 2 BUF2 $T=902100 769560 1 0 $X=902100 $Y=764140
X2989 3152 3279 1 2 BUF2 $T=903960 759480 1 0 $X=903960 $Y=754060
X2990 3341 3277 1 2 BUF2 $T=919460 779640 1 0 $X=919460 $Y=774220
X2991 3279 3512 1 2 BUF2 $T=944260 759480 1 0 $X=944260 $Y=754060
X2992 3603 3646 1 2 BUF2 $T=987040 809880 0 0 $X=987040 $Y=809500
X2993 3678 565 1 2 BUF2 $T=1016180 719160 0 0 $X=1016180 $Y=718780
X2994 3707 3680 1 2 BUF2 $T=1037260 759480 1 180 $X=1034160 $Y=759100
X2995 3696 3707 1 2 BUF2 $T=1045320 769560 0 180 $X=1042220 $Y=764140
X2996 2389 315 2380 2 318 2327 1 AO22 $T=735940 739320 0 180 $X=730980 $Y=733900
X2997 45 824 1 2 INV3 $T=388120 870360 0 0 $X=388120 $Y=869980
X2998 976 1025 1 2 INV3 $T=415400 759480 1 0 $X=415400 $Y=754060
X2999 47 135 1 2 INV3 $T=489180 759480 1 0 $X=489180 $Y=754060
X3000 1358 156 1 2 INV3 $T=511500 890520 0 0 $X=511500 $Y=890140
X3001 1457 1369 1 2 INV3 $T=520800 759480 0 180 $X=518320 $Y=754060
X3002 1646 1659 1 2 INV3 $T=565440 759480 0 0 $X=565440 $Y=759100
X3003 1840 177 1 2 INV3 $T=611320 739320 0 180 $X=608840 $Y=733900
X3004 291 283 1 2 INV3 $T=705560 719160 0 0 $X=705560 $Y=718780
X3005 2319 2355 1 2 INV3 $T=726020 749400 0 0 $X=726020 $Y=749020
X3006 2259 2383 1 2 INV3 $T=735940 809880 1 180 $X=733460 $Y=809500
X3007 2918 434 1 2 INV3 $T=857460 880440 1 0 $X=857460 $Y=875020
X3008 3025 3086 1 2 INV3 $T=871100 769560 0 0 $X=871100 $Y=769180
X3009 3051 442 1 2 INV3 $T=872960 880440 1 0 $X=872960 $Y=875020
X3010 3133 3179 1 2 INV3 $T=894040 779640 1 0 $X=894040 $Y=774220
X3011 3681 3662 1 2 INV3 $T=1018040 749400 1 0 $X=1018040 $Y=743980
X3012 991 937 1 2 BUF6 $T=415400 779640 1 180 $X=407960 $Y=779260
X3013 965 976 1 2 BUF6 $T=411060 749400 0 0 $X=411060 $Y=749020
X3014 56 965 1 2 BUF6 $T=411680 749400 1 0 $X=411680 $Y=743980
X3015 63 1039 1 2 BUF6 $T=417880 729240 0 0 $X=417880 $Y=728860
X3016 220 1837 1 2 BUF6 $T=626200 779640 0 0 $X=626200 $Y=779260
X3017 1980 2063 1 2 BUF6 $T=653480 769560 1 0 $X=653480 $Y=764140
X3018 2437 351 1 2 BUF6 $T=760740 860280 1 0 $X=760740 $Y=854860
X3019 417 2935 1 2 BUF6 $T=843200 880440 0 0 $X=843200 $Y=880060
X3020 3350 3170 1 2 BUF6 $T=920700 789720 0 0 $X=920700 $Y=789340
X3021 3679 3699 1 2 BUF6 $T=1026720 809880 1 0 $X=1026720 $Y=804460
X3022 565 567 1 2 BUF6 $T=1035400 719160 1 180 $X=1027960 $Y=718780
X3023 3697 3696 1 2 BUF6 $T=1037260 789720 1 0 $X=1037260 $Y=784300
X3024 3699 3697 1 2 BUF6 $T=1044700 799800 0 180 $X=1037260 $Y=794380
X3025 806 1 30 799 764 785 2 OAI22S $T=370760 759480 1 180 $X=367040 $Y=759100
X3026 798 1 30 785 733 806 2 OAI22S $T=367660 769560 1 0 $X=367660 $Y=764140
X3027 801 1 30 31 781 818 2 OAI22S $T=368280 729240 1 0 $X=368280 $Y=723820
X3028 837 1 857 850 770 846 2 OAI22S $T=383160 769560 1 180 $X=379440 $Y=769180
X3029 843 1 850 855 832 837 2 OAI22S $T=383160 789720 1 180 $X=379440 $Y=789340
X3030 930 1 933 937 744 963 2 OAI22S $T=399900 759480 0 0 $X=399900 $Y=759100
X3031 1018 1 1012 937 1002 993 2 OAI22S $T=413540 769560 0 180 $X=409820 $Y=764140
X3032 1015 1 1013 994 952 991 2 OAI22S $T=413540 799800 0 180 $X=409820 $Y=794380
X3033 1015 1 1003 1021 1022 991 2 OAI22S $T=411680 799800 0 0 $X=411680 $Y=799420
X3034 1015 1 994 1020 962 991 2 OAI22S $T=416020 789720 1 180 $X=412300 $Y=789340
X3035 955 1 1099 1108 1056 1093 2 OAI22S $T=434620 759480 0 0 $X=434620 $Y=759100
X3036 297 1 295 287 2288 2257 2 OAI22S $T=714860 729240 0 180 $X=711140 $Y=723820
X3037 2257 1 295 287 2297 2301 2 OAI22S $T=711140 729240 0 0 $X=711140 $Y=728860
X3038 2377 1 332 2403 2414 2422 2 OAI22S $T=740280 749400 0 0 $X=740280 $Y=749020
X3039 2336 1 332 2403 2461 2459 2 OAI22S $T=747100 769560 1 0 $X=747100 $Y=764140
X3040 2450 1 332 336 2469 2377 2 OAI22S $T=755160 729240 0 180 $X=751440 $Y=723820
X3041 3089 1 3033 450 3148 3127 2 OAI22S $T=886600 890520 0 180 $X=882880 $Y=885100
X3042 3133 1 3204 3210 3216 3179 2 OAI22S $T=892800 789720 1 0 $X=892800 $Y=784300
X3043 3186 1 3048 3197 3220 3083 2 OAI22S $T=895900 749400 1 0 $X=895900 $Y=743980
X3044 3178 1 3033 470 3225 3202 2 OAI22S $T=899620 890520 1 180 $X=895900 $Y=890140
X3045 3257 1 3195 3200 474 3197 2 OAI22S $T=900860 739320 1 180 $X=897140 $Y=738940
X3046 3296 1 3271 3277 3287 3289 2 OAI22S $T=910780 769560 1 180 $X=907060 $Y=769180
X3047 3373 1 3195 3200 3352 3349 2 OAI22S $T=921940 739320 1 180 $X=918220 $Y=738940
X3048 3271 1 3443 3435 3465 3471 2 OAI22S $T=935580 779640 1 0 $X=935580 $Y=774220
X3049 3525 1 3341 3511 3513 3472 2 OAI22S $T=949840 799800 0 180 $X=946120 $Y=794380
X3050 3530 1 3195 3521 523 3505 2 OAI22S $T=951080 739320 0 180 $X=947360 $Y=733900
X3051 3511 1 3524 3435 3519 3495 2 OAI22S $T=951080 789720 0 180 $X=947360 $Y=784300
X3052 3511 1 3533 3435 3545 3549 2 OAI22S $T=951080 779640 0 0 $X=951080 $Y=779260
X3053 3547 1 3195 3521 3544 3530 2 OAI22S $T=956660 739320 0 180 $X=952940 $Y=733900
X3054 817 2 898 979 952 1 730 FA1S $T=404240 799800 0 180 $X=392460 $Y=794380
X3055 2758 2 2748 2765 2745 1 2797 FA1S $T=810960 779640 1 0 $X=810960 $Y=774220
X3056 2780 2 2856 2849 2783 1 2781 FA1S $T=832040 759480 1 180 $X=820260 $Y=759100
X3057 412 2 2888 2843 2743 1 2790 FA1S $T=840100 739320 0 180 $X=828320 $Y=733900
X3058 408 2 2887 2848 2770 1 420 FA1S $T=829560 729240 1 0 $X=829560 $Y=723820
X3059 3564 2 3584 3427 3513 1 3596 FA1S $T=954180 799800 0 0 $X=954180 $Y=799420
X3060 937 996 1 2 INV4 $T=411060 759480 1 0 $X=411060 $Y=754060
X3061 193 190 1 2 INV4 $T=587140 739320 0 180 $X=584040 $Y=733900
X3062 190 1358 1 2 INV4 $T=585900 739320 0 0 $X=585900 $Y=738940
X3063 1886 209 1 2 INV4 $T=617520 759480 0 180 $X=614420 $Y=754060
X3064 2383 2437 1 2 INV4 $T=756400 809880 0 0 $X=756400 $Y=809500
X3065 210 2635 1 2 INV4 $T=782440 840120 0 0 $X=782440 $Y=839740
X3066 2673 373 1 2 INV4 $T=792360 809880 0 0 $X=792360 $Y=809500
X3067 3580 3578 1 2 INV4 $T=962240 890520 1 180 $X=959140 $Y=890140
X3068 549 3603 1 2 INV4 $T=969060 809880 1 180 $X=965960 $Y=809500
X3069 603 599 1 596 2 OR2T $T=318680 759480 0 180 $X=312480 $Y=754060
X3070 635 636 1 624 2 OR2T $T=331080 739320 0 180 $X=324880 $Y=733900
X3071 2679 2650 1 2738 2 OR2T $T=802900 739320 1 0 $X=802900 $Y=733900
X3072 3066 3054 1 3026 2 OR2T $T=869860 850200 0 180 $X=863660 $Y=844780
X3073 3613 3624 1 553 2 OR2T $T=972780 719160 0 0 $X=972780 $Y=718780
X3074 3632 3620 1 555 2 OR2T $T=976500 729240 0 0 $X=976500 $Y=728860
X3075 58 989 986 960 2 55 1 AOI13HS $T=411060 729240 0 180 $X=407340 $Y=723820
X3076 2235 2338 2334 2331 2 2319 1 AOI13HS $T=723540 729240 1 180 $X=719820 $Y=728860
X3077 3117 3235 3249 3232 2 3179 1 AOI13HS $T=902100 779640 1 180 $X=898380 $Y=779260
X3078 610 603 602 1 2 600 OA12 $T=316820 749400 1 180 $X=313100 $Y=749020
X3079 2387 2403 2410 1 2 2424 OA12 $T=738420 779640 1 0 $X=738420 $Y=774220
X3080 2403 2355 2442 1 2 2454 OA12 $T=745240 759480 0 0 $X=745240 $Y=759100
X3081 2560 2540 2526 1 2 2527 OA12 $T=769420 769560 1 180 $X=765700 $Y=769180
X3082 2690 2669 2630 1 2 2704 OA12 $T=796080 769560 1 0 $X=796080 $Y=764140
X3083 2762 2766 2772 1 2 2776 OA12 $T=817160 860280 1 0 $X=817160 $Y=854860
X3084 2985 2940 2958 1 2 2890 OA12 $T=854980 850200 1 180 $X=851260 $Y=849820
X3085 2964 2936 2950 1 2 2916 OA12 $T=858700 759480 1 180 $X=854980 $Y=759100
X3086 3011 2994 3017 1 2 3010 OA12 $T=861180 729240 1 0 $X=861180 $Y=723820
X3087 3133 3048 3137 1 2 2980 OA12 $T=884120 769560 1 180 $X=880400 $Y=769180
X3088 3270 470 3328 1 2 3342 OA12 $T=911400 890520 0 0 $X=911400 $Y=890140
X3089 934 933 1 917 788 911 2 OAI22H $T=399280 739320 1 180 $X=391840 $Y=738940
X3090 925 933 1 934 797 917 2 OAI22H $T=400520 749400 0 180 $X=393080 $Y=743980
X3091 911 933 1 945 826 939 2 OAI22H $T=394940 739320 1 0 $X=394940 $Y=733900
X3092 933 939 1 945 52 958 2 OAI22H $T=396180 729240 0 0 $X=396180 $Y=728860
X3093 3271 3395 1 3277 511 3423 2 OAI22H $T=923800 769560 1 0 $X=923800 $Y=764140
X3094 2841 2687 2884 417 1 2 QDFFRBP $T=829560 840120 1 0 $X=829560 $Y=834700
X3095 2975 2687 2914 424 1 2 QDFFRBP $T=856220 840120 0 180 $X=843820 $Y=834700
X3096 2921 360 2902 3001 1 2 QDFFRBP $T=847540 789720 1 0 $X=847540 $Y=784300
X3097 2860 360 2902 3025 1 2 QDFFRBP $T=850640 779640 0 0 $X=850640 $Y=779260
X3098 3070 2687 3084 3111 1 2 QDFFRBP $T=872960 830040 0 0 $X=872960 $Y=829660
X3099 2850 2687 3106 3174 1 2 QDFFRBP $T=876060 789720 0 0 $X=876060 $Y=789340
X3100 2632 360 2729 2 1 2744 QDFFRBS $T=797320 789720 1 0 $X=797320 $Y=784300
X3101 1265 1270 1 1278 1281 2 1258 1204 1279 OAI222S $T=476780 749400 1 0 $X=476780 $Y=743980
X3102 1265 1297 1 1276 1281 2 116 1200 1279 OAI222S $T=484840 739320 1 180 $X=479260 $Y=738940
X3103 1265 1318 1 126 1281 2 124 1256 1279 OAI222S $T=485460 749400 1 0 $X=485460 $Y=743980
X3104 1336 1335 1 1313 1325 2 1260 1136 1322 OAI222S $T=492900 789720 0 180 $X=487320 $Y=784300
X3105 1336 1300 1 1343 1325 2 1288 1161 1322 OAI222S $T=490420 779640 1 0 $X=490420 $Y=774220
X3106 1336 1329 1 1359 1325 2 1305 1106 1322 OAI222S $T=500340 789720 0 180 $X=494760 $Y=784300
X3107 1369 1393 1 144 1382 2 138 1264 1374 OAI222S $T=506540 739320 0 180 $X=500960 $Y=733900
X3108 1336 1413 1 1412 1325 2 1401 1170 1435 OAI222S $T=509640 769560 0 0 $X=509640 $Y=769180
X3109 1369 150 1 151 1382 2 147 1255 1374 OAI222S $T=510260 739320 1 0 $X=510260 $Y=733900
X3110 1336 1455 1 157 1325 2 1426 1165 1435 OAI222S $T=522040 769560 0 180 $X=516460 $Y=764140
X3111 1369 1437 1 161 1382 2 159 1248 1374 OAI222S $T=518320 739320 1 0 $X=518320 $Y=733900
X3112 1336 1476 1 1470 1325 2 1438 1171 1435 OAI222S $T=526380 769560 1 180 $X=520800 $Y=769180
X3113 1504 167 1 165 1382 2 164 1199 1374 OAI222S $T=533820 739320 0 180 $X=528240 $Y=733900
X3114 1369 1528 1 1535 1540 2 1510 1164 1435 OAI222S $T=536300 759480 0 0 $X=536300 $Y=759100
X3115 1369 1529 1 1536 1540 2 1543 1205 1435 OAI222S $T=536300 769560 1 0 $X=536300 $Y=764140
X3116 1567 1322 1 1540 1586 2 1594 1104 1589 OAI222S $T=555520 799800 0 180 $X=549940 $Y=794380
X3117 1658 1504 1 1641 1682 2 1679 181 1653 OAI222S $T=567300 739320 1 0 $X=567300 $Y=733900
X3118 1504 1679 1 1658 1682 2 1691 187 1653 OAI222S $T=576600 739320 1 0 $X=576600 $Y=733900
X3119 1504 1847 1 1797 1682 2 1794 204 1653 OAI222S $T=612560 739320 1 180 $X=606980 $Y=738940
X3120 1913 1894 1 1837 1824 2 1887 213 1589 OAI222S $T=626820 789720 0 180 $X=621240 $Y=784300
X3121 1589 2177 1 1729 2171 2 2066 2176 1894 OAI222S $T=686340 799800 0 180 $X=680760 $Y=794380
X3122 2150 2200 1 2171 1765 2 2126 2204 1589 OAI222S $T=689440 799800 1 0 $X=689440 $Y=794380
X3123 282 2035 1 1719 2236 2 2178 2217 2200 OAI222S $T=696880 850200 1 0 $X=696880 $Y=844780
X3124 2234 2112 1 1712 2171 2 2175 2249 2259 OAI222S $T=698740 809880 1 0 $X=698740 $Y=804460
X3125 1589 2047 1 1761 2171 2 2224 2250 2200 OAI222S $T=704940 799800 0 180 $X=699360 $Y=794380
X3126 2234 2079 1 1795 2171 2 2144 2238 2200 OAI222S $T=704940 809880 1 180 $X=699360 $Y=809500
X3127 282 2051 1 1714 2236 2 2183 2248 292 OAI222S $T=701840 850200 0 0 $X=701840 $Y=849820
X3128 282 2278 1 2294 2236 2 2231 2293 292 OAI222S $T=713000 850200 0 0 $X=713000 $Y=849820
X3129 282 2308 1 2268 301 2 2307 2315 292 OAI222S $T=714240 860280 0 0 $X=714240 $Y=859900
X3130 2265 2161 1 2318 2344 2 2345 2332 2259 OAI222S $T=719820 799800 0 0 $X=719820 $Y=799420
X3131 2265 2299 1 2230 2344 2 2186 2357 2259 OAI222S $T=726020 799800 0 0 $X=726020 $Y=799420
X3132 2265 2214 1 2273 2344 2 2350 2340 2259 OAI222S $T=726640 809880 0 0 $X=726640 $Y=809500
X3133 2265 2306 1 2292 2344 2 2264 2388 2397 OAI222S $T=730980 819960 1 0 $X=730980 $Y=814540
X3134 2265 2220 1 2289 2344 2 2269 2381 2259 OAI222S $T=731600 799800 0 0 $X=731600 $Y=799420
X3135 2500 2379 1 2405 2506 2 2444 2498 2437 OAI222S $T=761980 840120 1 180 $X=756400 $Y=839740
X3136 2500 2491 1 2463 2506 2 2464 2499 2437 OAI222S $T=761980 850200 1 180 $X=756400 $Y=849820
X3137 2500 2351 1 2363 2506 2 2409 2519 2437 OAI222S $T=756400 860280 0 0 $X=756400 $Y=859900
X3138 2500 2399 1 2348 2506 2 2359 2524 2437 OAI222S $T=766940 850200 0 180 $X=761360 $Y=844780
X3139 2558 354 1 340 301 2 2512 353 351 OAI222S $T=768800 900600 0 180 $X=763220 $Y=895180
X3140 2558 350 1 2438 301 2 2492 2541 351 OAI222S $T=770040 890520 1 180 $X=764460 $Y=890140
X3141 2558 2525 1 356 2506 2 339 2567 351 OAI222S $T=773760 870360 1 180 $X=768180 $Y=869980
X3142 2620 2483 1 2426 2621 2 2415 2636 2569 OAI222S $T=779960 809880 0 0 $X=779960 $Y=809500
X3143 2620 2443 1 2504 2621 2 2548 2632 2569 OAI222S $T=780580 809880 1 0 $X=780580 $Y=804460
X3144 2635 2570 1 2591 2621 2 2593 2625 351 OAI222S $T=786780 860280 0 180 $X=781200 $Y=854860
X3145 2635 2626 1 2600 2621 2 2634 2665 2660 OAI222S $T=784300 819960 0 0 $X=784300 $Y=819580
X3146 2635 2530 1 2607 2621 2 2497 2667 2660 OAI222S $T=795460 830040 0 180 $X=789880 $Y=824620
X3147 373 2604 1 2629 2661 2 2672 2689 2660 OAI222S $T=799180 809880 0 180 $X=793600 $Y=804460
X3148 373 2544 1 2595 376 2 2436 2691 2660 OAI222S $T=801660 799800 1 180 $X=796080 $Y=799420
X3149 2635 2686 1 2694 2661 2 2711 2724 2660 OAI222S $T=797320 819960 0 0 $X=797320 $Y=819580
X3150 2635 2708 1 2705 2661 2 2717 2719 2660 OAI222S $T=798560 819960 1 0 $X=798560 $Y=814540
X3151 82 78 87 2 1 93 94 78 87 102 589 ICV_12 $T=435860 900600 1 0 $X=435860 $Y=895180
X3152 1326 882 1337 2 1 1370 1373 882 1395 1403 589 ICV_12 $T=488560 830040 0 0 $X=488560 $Y=829660
X3153 1312 1339 1360 2 1 1376 1387 1339 1360 1427 589 ICV_12 $T=490420 779640 0 0 $X=490420 $Y=779260
X3154 1332 133 1367 2 1 1366 1390 133 1367 1431 589 ICV_12 $T=491040 749400 1 0 $X=491040 $Y=743980
X3155 1353 130 1315 2 1 1398 1400 130 1315 1451 589 ICV_12 $T=494760 880440 0 0 $X=494760 $Y=880060
X3156 1491 1339 1527 2 1 1538 1544 1339 1527 1592 589 ICV_12 $T=527620 789720 1 0 $X=527620 $Y=784300
X3157 1583 130 1609 2 1 1607 1623 130 1609 1678 589 ICV_12 $T=546840 880440 0 0 $X=546840 $Y=880060
X3158 1596 1339 1527 2 1 1625 1649 1339 1680 1700 589 ICV_12 $T=551180 789720 1 0 $X=551180 $Y=784300
X3159 1704 1339 1680 2 1 1746 1760 1339 1781 1785 589 ICV_12 $T=575360 789720 1 0 $X=575360 $Y=784300
X3160 1736 130 185 2 1 1774 1783 130 1751 1809 589 ICV_12 $T=581560 890520 1 0 $X=581560 $Y=885100
X3161 1769 1733 1798 2 1 1813 1822 1733 1798 1854 589 ICV_12 $T=590240 759480 1 0 $X=590240 $Y=754060
X3162 1915 198 1952 2 1 1893 1975 198 1952 2021 589 ICV_12 $T=625580 880440 0 0 $X=625580 $Y=880060
X3163 1949 1733 1979 2 1 1991 1998 1733 1979 2032 589 ICV_12 $T=630540 759480 1 0 $X=630540 $Y=754060
X3164 2036 1733 2085 2 1 2099 2102 1733 2085 2149 589 ICV_12 $T=655340 819960 0 0 $X=655340 $Y=819580
X3165 2169 2127 2147 2 1 2203 2217 2127 2147 290 589 ICV_12 $T=682000 769560 1 0 $X=682000 $Y=764140
X3166 2285 270 2247 2 1 2321 2343 270 308 2364 589 ICV_12 $T=710520 880440 1 0 $X=710520 $Y=875020
X3167 2353 270 2354 2 1 2413 2419 270 338 2472 589 ICV_12 $T=729740 870360 0 0 $X=729740 $Y=869980
X3168 2534 270 2583 2 1 2596 2598 270 2583 2645 589 ICV_12 $T=763220 880440 1 0 $X=763220 $Y=875020
X3169 2531 360 2728 2 1 2742 2731 360 2728 395 589 ICV_12 $T=796700 749400 0 0 $X=796700 $Y=749020
X3170 2676 2687 2749 2 1 2725 2665 2687 2755 2821 589 ICV_12 $T=803520 819960 0 0 $X=803520 $Y=819580
X3171 2746 360 2729 2 1 397 2774 360 2825 2848 589 ICV_12 $T=809100 789720 1 0 $X=809100 $Y=784300
X3172 2689 2687 2749 2 1 2816 2822 2687 2749 2857 589 ICV_12 $T=814680 809880 0 0 $X=814680 $Y=809500
X3173 2802 360 2732 2 1 2867 2867 360 2902 2920 589 ICV_12 $T=822740 769560 0 0 $X=822740 $Y=769180
X3174 1025 2 1 978 BUF3 $T=416020 769560 1 0 $X=416020 $Y=764140
X3175 2012 2 1 1980 BUF3 $T=645420 799800 1 0 $X=645420 $Y=794380
X3176 1943 2 1 2200 BUF3 $T=688200 789720 0 0 $X=688200 $Y=789340
X3177 304 2 1 2319 BUF3 $T=722920 719160 1 180 $X=719200 $Y=718780
X3178 47 50 1 2 INV6 $T=389980 759480 0 0 $X=389980 $Y=759100
X3179 964 27 935 2 1 1009 1028 27 935 1069 589 ICV_14 $T=403000 870360 0 0 $X=403000 $Y=869980
X3180 1553 133 1537 2 1 1608 1617 133 176 1665 589 ICV_14 $T=543740 729240 0 0 $X=543740 $Y=728860
X3181 1556 133 176 2 1 1590 1619 133 179 1670 589 ICV_14 $T=544360 719160 0 0 $X=544360 $Y=718780
X3182 1666 1339 1632 2 1 1716 1717 1339 1632 1756 589 ICV_14 $T=567300 819960 0 0 $X=567300 $Y=819580
X3183 1667 130 1660 2 1 1720 1698 130 1660 1771 589 ICV_14 $T=567300 850200 1 0 $X=567300 $Y=844780
X3184 1744 1339 1750 2 1 1782 1791 1339 1772 1845 589 ICV_14 $T=583420 830040 0 0 $X=583420 $Y=829660
X3185 1743 1339 1750 2 1 1800 1810 1733 1762 1844 589 ICV_14 $T=587140 819960 1 0 $X=587140 $Y=814540
X3186 1811 198 1842 2 1 1860 1869 198 1842 1900 589 ICV_14 $T=599540 850200 0 0 $X=599540 $Y=849820
X3187 2010 198 1982 2 1 2052 2059 198 2050 2091 589 ICV_14 $T=644800 830040 0 0 $X=644800 $Y=829660
X3188 2017 198 2050 2 1 2061 2068 198 2050 2086 589 ICV_14 $T=647280 850200 1 0 $X=647280 $Y=844780
X3189 2062 1733 2098 2 1 2111 2118 1733 2098 2163 589 ICV_14 $T=658440 789720 1 0 $X=658440 $Y=784300
X3190 2322 270 2354 2 1 2366 2376 270 2354 2420 589 ICV_14 $T=718580 860280 1 0 $X=718580 $Y=854860
X3191 2369 2127 2391 2 1 2412 2421 2127 2391 2476 589 ICV_14 $T=729740 840120 0 0 $X=729740 $Y=839740
X3192 2524 360 2729 2 1 2741 2667 360 2729 2792 589 ICV_14 $T=796700 779640 0 0 $X=796700 $Y=779260
X3193 2971 2687 2851 2 1 440 3055 2687 3063 3080 589 ICV_14 $T=854360 819960 1 0 $X=854360 $Y=814540
X3194 3201 2687 3221 2 1 3331 3102 2687 3221 3383 589 ICV_14 $T=903340 809880 0 0 $X=903340 $Y=809500
X3195 3272 1 3527 2 BUF4CK $T=946120 759480 0 0 $X=946120 $Y=759100
X3196 2063 2147 1 2 BUF4 $T=673940 769560 1 0 $X=673940 $Y=764140
X3197 3646 3679 1 2 BUF4 $T=1023000 799800 0 0 $X=1023000 $Y=799420
X3198 747 757 731 2 1 728 XOR3 $T=361460 739320 0 180 $X=350300 $Y=733900
X3199 781 794 776 2 1 24 XOR3 $T=373860 719160 1 180 $X=362700 $Y=718780
X3200 3434 3417 3431 2 1 3475 XOR3 $T=932480 880440 0 0 $X=932480 $Y=880060
X3201 3612 3609 3601 2 1 3613 XOR3 $T=970920 739320 0 0 $X=970920 $Y=738940
X3202 621 607 619 615 1 2 ND3P $T=323020 799800 0 180 $X=318060 $Y=794380
X3203 667 690 670 685 1 2 ND3P $T=333560 789720 0 0 $X=333560 $Y=789340
X3204 2656 2649 2647 2651 1 2 ND3P $T=791740 759480 1 180 $X=786780 $Y=759100
X3205 2735 2722 2658 2738 1 2 ND3P $T=808480 739320 1 180 $X=803520 $Y=738940
X3206 2812 2793 2787 2799 1 2 ND3P $T=827080 850200 0 180 $X=822120 $Y=844780
X3207 3020 446 445 3053 1 2 ND3P $T=864280 719160 0 0 $X=864280 $Y=718780
X3208 3537 3528 3553 534 1 2 ND3P $T=954800 880440 0 180 $X=949840 $Y=875020
X3209 3414 3593 3575 3554 1 2 ND3P $T=958520 870360 1 0 $X=958520 $Y=864940
X3210 3577 3592 3428 3554 1 2 ND3P $T=960380 850200 0 0 $X=960380 $Y=849820
X3211 3592 3429 3595 3582 1 2 ND3P $T=967200 860280 0 180 $X=962240 $Y=854860
X3212 3608 3627 3593 3625 1 2 ND3P $T=969060 870360 1 0 $X=969060 $Y=864940
X3213 684 677 631 1 2 OR2P $T=337280 779640 0 180 $X=333560 $Y=774220
X3214 917 925 918 1 2 OR2P $T=396800 749400 1 180 $X=393080 $Y=749020
X3215 2523 2502 2614 1 2 OR2P $T=773760 779640 1 0 $X=773760 $Y=774220
X3216 2996 2923 3007 1 2 OR2P $T=858700 850200 1 0 $X=858700 $Y=844780
X3217 545 546 3611 1 2 OR2P $T=965340 900600 1 0 $X=965340 $Y=895180
X3218 3574 2 1 3611 3577 NR2F $T=963480 890520 1 0 $X=963480 $Y=885100
X3219 630 6 5 10 3747 1 2 DFFRBP $T=324880 719160 1 180 $X=310620 $Y=718780
X3220 3440 2687 3425 3748 508 1 2 DFFRBP $T=940540 819960 1 180 $X=926280 $Y=819580
X3221 3604 2687 3420 538 3749 1 2 DFFRBP $T=968440 830040 0 180 $X=954180 $Y=824620
X3222 3619 2687 3603 543 3750 1 2 DFFRBP $T=975880 819960 0 180 $X=961620 $Y=814540
X3223 1213 1 2 1238 INV3CK $T=466860 850200 0 0 $X=466860 $Y=849820
X3224 1382 1 2 129 INV3CK $T=502200 739320 0 0 $X=502200 $Y=738940
X3225 3569 1 2 3574 INV3CK $T=959760 880440 0 0 $X=959760 $Y=880060
X3226 549 541 1 2 INV12 $T=963480 809880 1 180 $X=956040 $Y=809500
X3227 537 534 1 539 3580 2 OAI12HP $T=952940 900600 1 0 $X=952940 $Y=895180
X3228 3483 3497 1 3510 3506 3504 2 OAI112HS $T=949840 850200 0 180 $X=945500 $Y=844780
X3229 3534 2687 3420 531 1 2 3751 DFFRBN $T=957900 819960 1 180 $X=944880 $Y=819580
X3230 3538 2687 3420 532 1 2 3752 DFFRBN $T=958520 830040 1 180 $X=945500 $Y=829660
X3231 2712 1 2730 2722 2 381 ND3HT $T=809720 729240 1 180 $X=802280 $Y=728860
X3232 3007 1 3026 2823 2 3038 ND3HT $T=868620 840120 0 180 $X=861180 $Y=834700
X3233 3081 1 3046 3038 2 3114 ND3HT $T=881020 840120 0 180 $X=873580 $Y=834700
X3234 3293 1 3114 3303 2 3318 ND3HT $T=915120 840120 0 180 $X=907680 $Y=834700
X3235 3401 1 3392 3318 2 3414 ND3HT $T=932480 840120 0 180 $X=925040 $Y=834700
X3236 3401 1 3392 3318 2 3428 ND3HT $T=934960 840120 1 180 $X=927520 $Y=839740
X3237 3523 1 3517 3492 2 3526 ND3HT $T=952320 870360 0 180 $X=944880 $Y=864940
X3238 862 864 767 844 1 37 2 AOI22S $T=387500 739320 1 180 $X=383780 $Y=738940
X3239 1044 1050 68 1052 1 1062 2 AOI22S $T=420360 739320 0 0 $X=420360 $Y=738940
X3240 1079 1052 810 1059 1 1062 2 AOI22S $T=427800 739320 1 180 $X=424080 $Y=738940
X3241 1083 1079 787 1052 1 1062 2 AOI22S $T=431520 749400 0 180 $X=427800 $Y=743980
X3242 1072 1075 904 1078 1 1082 2 AOI22S $T=427800 759480 0 0 $X=427800 $Y=759100
X3243 1086 1075 769 1076 1 1072 2 AOI22S $T=431520 769560 0 180 $X=427800 $Y=764140
X3244 1078 1075 772 1083 1 1072 2 AOI22S $T=429040 759480 1 0 $X=429040 $Y=754060
X3245 1076 1082 740 1075 1 1072 2 AOI22S $T=433380 769560 1 0 $X=433380 $Y=764140
X3246 1062 1114 83 1125 1 1092 2 AOI22S $T=436480 729240 0 0 $X=436480 $Y=728860
X3247 1183 1114 101 1191 1 99 2 AOI22S $T=455700 729240 1 0 $X=455700 $Y=723820
X3248 99 1114 1206 75 1 1224 2 AOI22S $T=461280 729240 1 0 $X=461280 $Y=723820
X3249 2393 2471 2432 2360 1 2465 2 AOI22S $T=754540 759480 1 180 $X=750820 $Y=759100
X3250 2402 2467 2529 2471 1 2465 2 AOI22S $T=761360 749400 1 180 $X=757640 $Y=749020
X3251 2416 2471 2536 2441 1 2465 2 AOI22S $T=765080 759480 1 180 $X=761360 $Y=759100
X3252 2520 2470 2538 2528 1 2516 2 AOI22S $T=764460 729240 0 0 $X=764460 $Y=728860
X3253 2470 2439 2539 2528 1 2516 2 AOI22S $T=764460 739320 1 0 $X=764460 $Y=733900
X3254 355 2549 2562 2520 1 344 2 AOI22S $T=768800 729240 0 180 $X=765080 $Y=723820
X3255 428 2938 2946 2900 1 2932 2 AOI22S $T=851880 860280 1 180 $X=848160 $Y=859900
X3256 2941 2938 2895 2953 1 2932 2 AOI22S $T=850020 870360 1 0 $X=850020 $Y=864940
X3257 2997 2988 2949 2976 1 3009 2 AOI22S $T=858700 870360 0 0 $X=858700 $Y=869980
X3258 3008 3018 2978 3015 1 2920 2 AOI22S $T=861800 759480 1 0 $X=861800 $Y=754060
X3259 3039 3047 2987 3018 1 2920 2 AOI22S $T=865520 769560 1 0 $X=865520 $Y=764140
X3260 3091 3068 3074 3018 1 3069 2 AOI22S $T=874200 749400 1 180 $X=870480 $Y=749020
X3261 3092 3060 3065 3079 1 3009 2 AOI22S $T=874200 870360 0 180 $X=870480 $Y=864940
X3262 3160 3092 3140 3079 1 3009 2 AOI22S $T=882260 870360 0 180 $X=878540 $Y=864940
X3263 3203 3079 3176 3160 1 3168 2 AOI22S $T=890320 870360 0 180 $X=886600 $Y=864940
X3264 3191 3169 3187 3132 1 3069 2 AOI22S $T=892800 749400 0 180 $X=889080 $Y=743980
X3265 473 3079 3219 3203 1 3168 2 AOI22S $T=895900 870360 0 180 $X=892180 $Y=864940
X3266 3283 3191 3258 3267 1 3069 2 AOI22S $T=906440 739320 1 180 $X=902720 $Y=738940
X3267 3313 3267 3292 3283 1 3307 2 AOI22S $T=913260 739320 0 180 $X=909540 $Y=733900
X3268 496 3147 3306 473 1 3168 2 AOI22S $T=916980 880440 1 180 $X=913260 $Y=880060
X3269 498 3147 3355 496 1 3168 2 AOI22S $T=919460 890520 0 180 $X=915740 $Y=885100
X3270 499 3147 3379 498 1 3168 2 AOI22S $T=920700 890520 1 180 $X=916980 $Y=890140
X3271 494 3147 3345 499 1 3168 2 AOI22S $T=917600 900600 1 0 $X=917600 $Y=895180
X3272 3267 3307 3381 3372 1 3313 2 AOI22S $T=923800 739320 0 180 $X=920080 $Y=733900
X3273 3424 3267 509 3372 1 3307 2 AOI22S $T=928760 739320 0 180 $X=925040 $Y=733900
X3274 3437 3424 3433 3267 1 3307 2 AOI22S $T=933720 739320 0 180 $X=930000 $Y=733900
X3275 3486 3468 3469 3437 1 3307 2 AOI22S $T=941160 739320 0 180 $X=937440 $Y=733900
X3276 3460 3468 526 3486 1 3307 2 AOI22S $T=946120 739320 0 180 $X=942400 $Y=733900
X3277 3354 3170 3301 3331 2 1 NR3H $T=918220 799800 1 180 $X=912640 $Y=799420
X3278 51 1 2 830 BUF1CK $T=400520 729240 0 180 $X=398040 $Y=723820
X3279 63 1 2 960 BUF1CK $T=417880 729240 1 180 $X=415400 $Y=728860
X3280 1374 1 2 1435 BUF1CK $T=516460 739320 0 0 $X=516460 $Y=738940
X3281 2247 1 2 2201 BUF1CK $T=703700 880440 0 0 $X=703700 $Y=880060
X3282 2900 1 2 430 BUF1CK $T=850640 900600 1 0 $X=850640 $Y=895180
X3283 3172 1 2 3015 BUF1CK $T=889700 769560 0 180 $X=887220 $Y=764140
X3284 2696 1 2 3198 BUF1CK $T=890940 779640 0 0 $X=890940 $Y=779260
X3285 3250 1 2 3162 BUF1CK $T=900860 789720 1 0 $X=900860 $Y=784300
X3286 2935 1 2 480 BUF8CK $T=896520 890520 1 0 $X=896520 $Y=885100
X3287 699 710 1 716 652 2 OAI12H $T=341620 749400 0 0 $X=341620 $Y=749020
X3288 2599 2547 1 2614 2669 2 OAI12H $T=779340 769560 0 0 $X=779340 $Y=769180
X3289 2868 2863 1 2853 2766 2 OAI12H $T=835760 850200 1 180 $X=829560 $Y=849820
X3290 2969 2929 1 2995 2994 2 OAI12H $T=855600 739320 1 0 $X=855600 $Y=733900
X3291 3195 3186 1 3177 3141 2 OAI12H $T=894040 749400 1 180 $X=887840 $Y=749020
X3292 3213 3223 1 3206 3242 2 OAI12H $T=894660 840120 0 0 $X=894660 $Y=839740
X3293 3205 3233 1 3251 3261 2 OAI12H $T=896520 830040 0 0 $X=896520 $Y=829660
X3294 3172 1 3001 3137 3075 2 ND3S $T=889080 779640 0 180 $X=886600 $Y=774220
X3295 936 918 2 789 904 1 AOI12H $T=398660 759480 0 180 $X=392460 $Y=754060
X3296 2456 2527 2 2547 2507 1 AOI12H $T=760740 779640 0 0 $X=760740 $Y=779260
X3297 2892 2890 2 2863 2879 1 AOI12H $T=841960 850200 1 180 $X=835760 $Y=849820
X3298 2854 2771 2806 1 2 2827 HA1 $T=835760 759480 0 180 $X=827700 $Y=754060
X3299 796 27 824 2 1 835 842 847 589 ICV_17 $T=367040 870360 0 0 $X=367040 $Y=869980
X3300 919 882 943 2 1 970 970 931 589 ICV_17 $T=393080 830040 1 0 $X=393080 $Y=824620
X3301 948 882 886 2 1 1006 1006 1014 589 ICV_17 $T=399280 850200 0 0 $X=399280 $Y=849820
X3302 1060 882 1029 2 1 1103 1103 1077 589 ICV_17 $T=423460 830040 1 0 $X=423460 $Y=824620
X3303 1135 882 1090 2 1 1176 1176 1128 589 ICV_17 $T=442060 830040 1 0 $X=442060 $Y=824620
X3304 1187 882 1154 2 1 1222 1222 1235 589 ICV_17 $T=456320 769560 1 0 $X=456320 $Y=764140
X3305 1245 882 1227 2 1 1302 1242 1259 589 ICV_17 $T=471820 809880 0 0 $X=471820 $Y=809500
X3306 1430 1339 1414 2 1 1415 1478 1477 589 ICV_17 $T=513360 809880 0 0 $X=513360 $Y=809500
X3307 1572 1339 1595 2 1 1615 1615 1599 589 ICV_17 $T=544980 830040 0 0 $X=544980 $Y=829660
X3308 1673 1339 1632 2 1 1726 1726 1714 589 ICV_17 $T=568540 819960 1 0 $X=568540 $Y=814540
X3309 1690 130 1660 2 1 1775 1775 1701 589 ICV_17 $T=579700 860280 1 0 $X=579700 $Y=854860
X3310 1748 192 1703 2 1 1806 1737 1711 589 ICV_17 $T=588380 729240 1 0 $X=588380 $Y=723820
X3311 1912 198 1951 2 1 1962 1962 1930 589 ICV_17 $T=623720 850200 0 0 $X=623720 $Y=849820
X3312 1937 1733 1863 2 1 1986 1986 236 589 ICV_17 $T=628060 749400 1 0 $X=628060 $Y=743980
X3313 1974 1733 2012 2 1 1984 2019 2042 589 ICV_17 $T=641700 799800 0 0 $X=641700 $Y=799420
X3314 246 198 2044 2 1 2087 2087 252 589 ICV_17 $T=652240 900600 1 0 $X=652240 $Y=895180
X3315 2046 198 2078 2 1 2093 2093 2095 589 ICV_17 $T=653480 870360 1 0 $X=653480 $Y=864940
X3316 2041 198 2044 2 1 2105 2105 2051 589 ICV_17 $T=656580 870360 0 0 $X=656580 $Y=869980
X3317 2056 198 2092 2 1 2106 2104 258 589 ICV_17 $T=656580 890520 0 0 $X=656580 $Y=890140
X3318 2122 1733 2156 2 1 2172 2172 2161 589 ICV_17 $T=671460 809880 1 0 $X=671460 $Y=804460
X3319 2157 198 2188 2 1 2202 2202 2175 589 ICV_17 $T=679520 850200 0 0 $X=679520 $Y=849820
X3320 2266 2127 2314 2 1 2349 2349 2273 589 ICV_17 $T=713620 809880 0 0 $X=713620 $Y=809500
X3321 2274 2127 2277 2 1 2356 2356 2292 589 ICV_17 $T=716100 789720 0 0 $X=716100 $Y=789340
X3322 2303 2127 2277 2 1 2367 2367 2318 589 ICV_17 $T=718580 799800 1 0 $X=718580 $Y=794380
X3323 2337 2127 2391 2 1 2406 2406 2348 589 ICV_17 $T=727260 850200 1 0 $X=727260 $Y=844780
X3324 319 270 331 2 1 2428 2428 328 589 ICV_17 $T=732840 900600 1 0 $X=732840 $Y=895180
X3325 2396 2127 2433 2 1 2449 2449 2415 589 ICV_17 $T=736560 809880 0 0 $X=736560 $Y=809500
X3326 2429 2127 2433 2 1 2513 2513 2443 589 ICV_17 $T=748340 809880 1 0 $X=748340 $Y=804460
X3327 2481 270 338 2 1 2537 2537 350 589 ICV_17 $T=753300 870360 0 0 $X=753300 $Y=869980
X3328 2554 2127 2563 2 1 2609 2609 2607 589 ICV_17 $T=766320 830040 0 0 $X=766320 $Y=829660
X3329 2561 2127 2479 2 1 2611 2611 2604 589 ICV_17 $T=766940 809880 1 0 $X=766940 $Y=804460
X3330 2575 2127 2601 2 1 2644 2623 2600 589 ICV_17 $T=774380 850200 1 0 $X=774380 $Y=844780
X3331 2659 270 2648 2 1 2721 2726 380 589 ICV_17 $T=791740 890520 1 0 $X=791740 $Y=885100
X3332 2701 2687 2749 2 1 2760 2760 2711 589 ICV_17 $T=804140 830040 1 0 $X=804140 $Y=824620
X3333 2718 2687 2747 2 1 2777 2777 2705 589 ICV_17 $T=808480 809880 1 0 $X=808480 $Y=804460
X3334 103 97 1194 1177 2 1 1177 1130 1167 1152 589 ICV_18 $T=455700 880440 1 180 $X=450120 $Y=880060
X3335 1351 1299 1320 1331 2 1 1327 1299 1291 1316 589 ICV_18 $T=490420 890520 0 180 $X=484840 $Y=885100
X3336 1565 1561 1553 1412 2 1 1535 163 1508 165 589 ICV_18 $T=540020 739320 0 180 $X=534440 $Y=733900
X3337 1692 1622 1674 1637 2 1 1657 1622 1636 1604 589 ICV_18 $T=567300 870360 1 180 $X=561720 $Y=869980
X3338 186 1647 183 1587 2 1 182 1647 180 1640 589 ICV_18 $T=574740 719160 1 180 $X=569160 $Y=718780
X3339 1731 1668 1717 1684 2 1 1696 1668 1666 1651 589 ICV_18 $T=576600 830040 1 180 $X=571020 $Y=829660
X3340 1735 1668 1723 1709 2 1 1709 1668 1698 1696 589 ICV_18 $T=577220 840120 0 180 $X=571640 $Y=834700
X3341 1830 1796 1811 1773 2 1 1803 1796 1793 1701 589 ICV_18 $T=600160 860280 0 180 $X=594580 $Y=854860
X3342 2047 2000 2036 2029 2 1 1990 2000 1993 2008 589 ICV_18 $T=649760 819960 1 180 $X=644180 $Y=819580
X3343 2294 2227 2279 1719 2 1 2268 2227 2255 1714 589 ICV_18 $T=708660 850200 0 180 $X=703080 $Y=844780
X3344 2318 2209 2303 1765 2 1 2289 2209 2252 1761 589 ICV_18 $T=713000 799800 0 180 $X=707420 $Y=794380
X3345 2443 2378 2429 2220 2 1 2415 2378 2396 2186 589 ICV_18 $T=742760 809880 0 180 $X=737180 $Y=804460
X3346 339 2435 2419 2409 2 1 2409 2435 2425 2307 589 ICV_18 $T=747100 870360 0 180 $X=741520 $Y=864940
X3347 2626 2553 2615 2483 2 1 2600 2553 2574 2426 589 ICV_18 $T=777480 819960 1 180 $X=771900 $Y=819580
X3348 2717 2680 2707 2436 2 1 2694 2680 2682 2607 589 ICV_18 $T=798560 830040 1 180 $X=792980 $Y=829660
X3349 388 2716 2736 2717 2 1 380 2716 2677 2705 589 ICV_18 $T=804140 880440 0 180 $X=798560 $Y=875020
X3350 389 2716 2740 2686 2 1 382 2716 2715 2604 589 ICV_18 $T=806000 870360 0 180 $X=800420 $Y=864940
X3351 631 1 675 650 2 ND2T $T=331700 789720 1 0 $X=331700 $Y=784300
X3352 215 1 220 1886 2 ND2T $T=623720 769560 1 0 $X=623720 $Y=764140
X3353 215 1 1837 1943 2 ND2T $T=628680 789720 1 180 $X=623720 $Y=789340
X3354 2678 1 2649 2735 2 ND2T $T=796700 749400 0 180 $X=791740 $Y=743980
X3355 337 359 361 2 1 2663 XNR3 $T=777480 719160 0 0 $X=777480 $Y=718780
X3356 614 607 8 595 1 2 MXL2H $T=318060 799800 0 180 $X=309380 $Y=794380
X3357 713 690 17 689 1 2 MXL2H $T=347200 789720 1 180 $X=338520 $Y=789340
X3358 904 905 692 871 1 2 MXL2H $T=392460 759480 0 180 $X=383780 $Y=754060
X3359 2222 283 287 2244 1 2 MXL2H $T=696880 729240 1 0 $X=696880 $Y=723820
X3360 2312 2355 305 2328 1 2 MXL2H $T=729740 759480 0 180 $X=721060 $Y=754060
X3361 2200 1 2259 2 BUF6CK $T=702460 799800 0 0 $X=702460 $Y=799420
X3362 249 277 1 2 INV6CK $T=690680 830040 0 180 $X=685100 $Y=824620
X3363 1062 1059 2 1052 69 1044 1 AOI22H $T=427180 749400 0 180 $X=419740 $Y=743980
X3364 61 1011 67 61 2 1 1034 MAOI1H $T=424700 719160 1 180 $X=417260 $Y=718780
X3365 1031 978 991 1065 1 2 MXL2HP $T=415400 779640 0 0 $X=415400 $Y=779260
X3366 915 1 2 46 BUF3CK $T=395560 769560 0 180 $X=391220 $Y=764140
X3367 717 700 692 1 2 XNR2H $T=347820 739320 1 180 $X=339140 $Y=738940
X3368 700 694 724 1 2 XNR2H $T=339760 739320 1 0 $X=339760 $Y=733900
X3369 742 727 721 1 2 XNR2H $T=357120 729240 0 180 $X=348440 $Y=723820
X3370 727 21 728 1 2 XNR2H $T=349060 719160 0 0 $X=349060 $Y=718780
X3371 624 622 610 608 1 2 OA12P $T=323020 739320 0 180 $X=318680 $Y=733900
X3372 602 599 594 617 1 2 OA12P $T=323020 759480 0 180 $X=318680 $Y=754060
X3373 633 628 626 615 1 2 OA12P $T=324880 799800 1 180 $X=320540 $Y=799420
X3374 635 622 642 644 1 2 OA12P $T=324880 729240 0 0 $X=324880 $Y=728860
X3375 646 691 681 628 1 2 OA12P $T=341000 779640 1 180 $X=336660 $Y=779260
X3376 20 18 19 16 1 2 OA12P $T=345340 719160 1 180 $X=341000 $Y=718780
X3377 596 610 1 617 620 2 OAI12HT $T=307520 759480 0 0 $X=307520 $Y=759100
X3378 591 6 5 4 1 2 3753 DFFRBS $T=306900 719160 1 180 $X=293880 $Y=718780
.ENDS
***************************************
.SUBCKT ICV_20 1 2 3 4 5 6 7 8 9 10 11
** N=11 EP=11 IP=14 FDC=0
X0 1 2 3 4 5 6 QDFFRBN $T=11780 0 0 180 $X=0 $Y=-5420
X1 7 8 9 4 5 10 QDFFRBN $T=0 0 0 0 $X=0 $Y=-380
.ENDS
***************************************
.SUBCKT MUX2S B S VCC A GND O
** N=7 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MUX2 B S VCC GND O A
** N=7 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AOI12HP B2 B1 VCC O A1 GND
** N=7 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AO12P B2 B1 A1 O GND VCC
** N=7 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MAO222P A1 B1 C1 O GND VCC
** N=7 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AN3 I1 I2 I3 VCC GND O
** N=7 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OAI222H C1 C2 GND B1 B2 A2 O A1 VCC
** N=10 EP=9 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MAOI1 B1 B2 A1 A2 VCC GND O
** N=8 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT BUF8 I O GND VCC
** N=5 EP=4 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT XNR2HP I2 O I1 GND VCC
** N=6 EP=5 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT INV2CK I O GND VCC
** N=5 EP=4 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ND2F I2 I1 VCC O GND
** N=6 EP=5 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_21 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140
+ 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160
+ 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180
+ 181 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200
+ 201 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220
+ 221 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240
+ 241 242 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 259 260
+ 261 262 263 264 265 266 267 268 269 270 271 272 273 274 275 276 277 278 279 280
+ 281 282 283 284 285 286 287 288 289 290 291 292 293 294 295 296 297 298 299 300
+ 301 302 303 304 305 306 307 308 309 310 311 312 313 314 315 316 317 318 319 320
+ 321 322 323 324 325 326 327 328 329 330 331 332 333 334 335 336 337 338 339 340
+ 341 342 343 344 345 346 347 348 349 350 351 352 353 354 355 356 357 358 359 360
+ 361 362 363 364 365 366 367 368 369 370 371 372 373 374 375 376 377 378 379 380
+ 381 382 383 384 385 386 387 388 389 390 391 392 393 394 395 396 397 398 399 400
+ 401 402 403 404 405 406 407 408 409 410 411 412 413 414 415 416 417 418 419 420
+ 421 422 423 424 425 426 427 428 429 430 431 432 433 434 435 436 437 438 439 440
+ 441 442 443 444 445 446 447 448 449 450 451 452 453 454 455 456 457 458 459 460
+ 461 462 463 464 465 466 467 468 469 470 471 472 473 474 475 476 477 478 479 480
+ 481 482 483 484 485 486 487 488 489 490 491 492 493 494 495 496 497 498 499 500
+ 501 502 503 504 505 506 507 508 509 510 511 512 513 514 515 516 517 518 519 520
+ 521 522 523 524 525 526 527 528 529 530 531 532 533 534 535 536 537 538 539 540
+ 541 542 543 544 545 546 547 548 549 550 551 552 553 554 555 556 557 558 559 560
+ 561 562 563 564 565 566 567 568 569 570 571 572 573 574 575 576 577 578 579 580
+ 581 582 583 584 585 586 587 588 589 590 591 592 593 594 595 596 597 598 599 600
+ 601 602 603 604 605 606 607 608 609 610 611 612 613 614 615 616 617 618 619 620
+ 621 622 623 624 625 626 627 628 629 630 631 632 633 634 635 636 637 638 639 640
+ 641 642 643 644 645 646 647 648 649 650 651 652 653 654 655 656 657 658 659 660
+ 661 662 663 675
** N=4659 EP=664 IP=25820 FDC=0
X0 1121 1 2 997 BUF1S $T=352780 638520 1 180 $X=350300 $Y=638140
X1 1273 1 2 61 BUF1S $T=377580 547800 1 0 $X=377580 $Y=542380
X2 377 1 2 2781 BUF1S $T=713620 709080 1 180 $X=711140 $Y=708700
X3 2710 1 2 2830 BUF1S $T=713620 699000 1 0 $X=713620 $Y=693580
X4 3757 1 2 3786 BUF1S $T=878540 638520 1 0 $X=878540 $Y=633100
X5 553 1 2 3917 BUF1S $T=908300 547800 0 180 $X=905820 $Y=542380
X6 3864 1 2 4022 BUF1S $T=910160 628440 0 0 $X=910160 $Y=628060
X7 628 1 2 4335 BUF1S $T=995720 618360 1 180 $X=993240 $Y=617980
X8 587 1 2 632 BUF1S $T=1005640 598200 1 0 $X=1005640 $Y=592780
X9 834 2 1 738 BUF1 $T=298840 567960 1 180 $X=296360 $Y=567580
X10 918 2 1 842 BUF1 $T=314960 638520 1 180 $X=312480 $Y=638140
X11 942 2 1 7 BUF1 $T=319300 699000 1 180 $X=316820 $Y=698620
X12 983 2 1 939 BUF1 $T=327980 648600 0 180 $X=325500 $Y=643180
X13 985 2 1 29 BUF1 $T=326740 567960 1 0 $X=326740 $Y=562540
X14 985 2 1 834 BUF1 $T=329220 567960 1 180 $X=326740 $Y=567580
X15 1018 2 1 871 BUF1 $T=332320 668760 1 0 $X=332320 $Y=663340
X16 1083 2 1 942 BUF1 $T=345340 699000 0 180 $X=342860 $Y=693580
X17 1147 2 1 1092 BUF1 $T=354640 648600 0 0 $X=354640 $Y=648220
X18 1247 2 1 918 BUF1 $T=365180 618360 1 180 $X=362700 $Y=617980
X19 971 2 1 1035 BUF1 $T=372000 578040 0 0 $X=372000 $Y=577660
X20 1291 2 1 1177 BUF1 $T=380060 658680 1 180 $X=377580 $Y=658300
X21 1306 2 1 1209 BUF1 $T=381920 668760 0 180 $X=379440 $Y=663340
X22 1329 2 1 1186 BUF1 $T=386880 658680 0 180 $X=384400 $Y=653260
X23 1083 2 1 1303 BUF1 $T=390600 688920 0 180 $X=388120 $Y=683500
X24 1394 2 1 70 BUF1 $T=399280 719160 0 180 $X=396800 $Y=713740
X25 1247 2 1 1443 BUF1 $T=406100 618360 1 0 $X=406100 $Y=612940
X26 1415 2 1 1434 BUF1 $T=407960 578040 0 0 $X=407960 $Y=577660
X27 1415 2 1 1481 BUF1 $T=412920 588120 1 0 $X=412920 $Y=582700
X28 1525 2 1 1419 BUF1 $T=425940 557880 0 180 $X=423460 $Y=552460
X29 1525 2 1 1412 BUF1 $T=425940 567960 1 180 $X=423460 $Y=567580
X30 1481 2 1 1549 BUF1 $T=429040 578040 0 0 $X=429040 $Y=577660
X31 111 2 1 88 BUF1 $T=429660 709080 0 0 $X=429660 $Y=708700
X32 1549 2 1 103 BUF1 $T=432760 557880 0 180 $X=430280 $Y=552460
X33 1549 2 1 1358 BUF1 $T=432140 567960 1 0 $X=432140 $Y=562540
X34 1481 2 1 1641 BUF1 $T=445160 588120 1 0 $X=445160 $Y=582700
X35 1641 2 1 1680 BUF1 $T=450740 598200 0 0 $X=450740 $Y=597820
X36 1641 2 1 1679 BUF1 $T=453840 578040 1 0 $X=453840 $Y=572620
X37 1684 2 1 1590 BUF1 $T=456940 547800 1 180 $X=454460 $Y=547420
X38 1699 2 1 1720 BUF1 $T=466240 638520 0 0 $X=466240 $Y=638140
X39 1764 2 1 1757 BUF1 $T=482360 688920 1 180 $X=479880 $Y=688540
X40 1880 2 1 1822 BUF1 $T=496000 678840 1 180 $X=493520 $Y=678460
X41 1902 2 1 1861 BUF1 $T=500960 588120 0 180 $X=498480 $Y=582700
X42 1893 2 1 1891 BUF1 $T=499100 618360 1 0 $X=499100 $Y=612940
X43 1946 2 1 1880 BUF1 $T=507780 678840 1 180 $X=505300 $Y=678460
X44 1934 2 1 1893 BUF1 $T=510260 608280 0 180 $X=507780 $Y=602860
X45 1893 2 1 1959 BUF1 $T=512120 628440 1 0 $X=512120 $Y=623020
X46 1940 2 1 1968 BUF1 $T=514600 699000 0 0 $X=514600 $Y=698620
X47 175 2 1 197 BUF1 $T=520180 719160 0 180 $X=517700 $Y=713740
X48 1934 2 1 1996 BUF1 $T=522040 608280 0 0 $X=522040 $Y=607900
X49 1938 2 1 2004 BUF1 $T=527000 567960 1 180 $X=524520 $Y=567580
X50 175 2 1 2007 BUF1 $T=524520 699000 0 0 $X=524520 $Y=698620
X51 2007 2 1 1986 BUF1 $T=527000 699000 0 0 $X=527000 $Y=698620
X52 1959 2 1 2028 BUF1 $T=528240 638520 0 0 $X=528240 $Y=638140
X53 2041 2 1 1954 BUF1 $T=533820 658680 0 180 $X=531340 $Y=653260
X54 1959 2 1 2041 BUF1 $T=532580 658680 0 0 $X=532580 $Y=658300
X55 1934 2 1 2051 BUF1 $T=533200 598200 0 0 $X=533200 $Y=597820
X56 2041 2 1 1946 BUF1 $T=533820 668760 0 0 $X=533820 $Y=668380
X57 2058 2 1 1931 BUF1 $T=535680 598200 0 0 $X=535680 $Y=597820
X58 2002 2 1 2088 BUF1 $T=540020 628440 1 0 $X=540020 $Y=623020
X59 1946 2 1 2090 BUF1 $T=540640 678840 1 0 $X=540640 $Y=673420
X60 2052 2 1 2009 BUF1 $T=546220 668760 1 180 $X=543740 $Y=668380
X61 2057 2 1 1942 BUF1 $T=544980 598200 1 0 $X=544980 $Y=592780
X62 2028 2 1 2125 BUF1 $T=551180 638520 0 0 $X=551180 $Y=638140
X63 2150 2 1 2081 BUF1 $T=561720 608280 1 180 $X=559240 $Y=607900
X64 2051 2 1 2150 BUF1 $T=562960 608280 0 180 $X=560480 $Y=602860
X65 243 2 1 255 BUF1 $T=560480 719160 1 0 $X=560480 $Y=713740
X66 2051 2 1 2174 BUF1 $T=564200 608280 1 0 $X=564200 $Y=602860
X67 2172 2 1 2108 BUF1 $T=567300 688920 1 180 $X=564820 $Y=688540
X68 2123 2 1 2164 BUF1 $T=572880 588120 0 180 $X=570400 $Y=582700
X69 255 2 1 261 BUF1 $T=571640 709080 0 0 $X=571640 $Y=708700
X70 2207 2 1 2186 BUF1 $T=575360 648600 0 180 $X=572880 $Y=643180
X71 255 2 1 2226 BUF1 $T=575360 699000 0 0 $X=575360 $Y=698620
X72 2186 2 1 2148 BUF1 $T=577840 628440 1 0 $X=577840 $Y=623020
X73 2172 2 1 2146 BUF1 $T=578460 668760 0 0 $X=578460 $Y=668380
X74 2226 2 1 2172 BUF1 $T=581560 688920 1 180 $X=579080 $Y=688540
X75 2258 2 1 2147 BUF1 $T=582800 557880 1 180 $X=580320 $Y=557500
X76 2148 2 1 2237 BUF1 $T=580940 608280 1 0 $X=580940 $Y=602860
X77 2123 2 1 2233 BUF1 $T=581560 578040 1 0 $X=581560 $Y=572620
X78 2258 2 1 2214 BUF1 $T=587760 557880 1 180 $X=585280 $Y=557500
X79 272 2 1 2235 BUF1 $T=585280 709080 0 0 $X=585280 $Y=708700
X80 2207 2 1 2266 BUF1 $T=587760 638520 1 0 $X=587760 $Y=633100
X81 2226 2 1 2261 BUF1 $T=589000 688920 0 0 $X=589000 $Y=688540
X82 264 2 1 2258 BUF1 $T=590240 547800 0 0 $X=590240 $Y=547420
X83 2150 2 1 2282 BUF1 $T=590860 618360 0 0 $X=590860 $Y=617980
X84 2207 2 1 2293 BUF1 $T=592100 648600 0 0 $X=592100 $Y=648220
X85 261 2 1 277 BUF1 $T=594580 719160 1 0 $X=594580 $Y=713740
X86 2306 2 1 2252 BUF1 $T=599540 648600 0 180 $X=597060 $Y=643180
X87 2258 2 1 2312 BUF1 $T=603880 557880 1 0 $X=603880 $Y=552460
X88 2235 2 1 2319 BUF1 $T=603880 709080 1 0 $X=603880 $Y=703660
X89 2298 2 1 2320 BUF1 $T=605120 578040 0 0 $X=605120 $Y=577660
X90 2261 2 1 2316 BUF1 $T=605740 678840 1 0 $X=605740 $Y=673420
X91 2266 2 1 2353 BUF1 $T=606980 638520 1 0 $X=606980 $Y=633100
X92 2319 2 1 2330 BUF1 $T=608840 699000 0 0 $X=608840 $Y=698620
X93 2298 2 1 2360 BUF1 $T=609460 588120 1 0 $X=609460 $Y=582700
X94 2360 2 1 280 BUF1 $T=613180 567960 0 180 $X=610700 $Y=562540
X95 2312 2 1 2376 BUF1 $T=612560 547800 0 0 $X=612560 $Y=547420
X96 2282 2 1 2387 BUF1 $T=613800 628440 1 0 $X=613800 $Y=623020
X97 2330 2 1 2364 BUF1 $T=614420 678840 0 0 $X=614420 $Y=678460
X98 277 2 1 296 BUF1 $T=615660 719160 1 0 $X=615660 $Y=713740
X99 2387 2 1 2306 BUF1 $T=619380 638520 0 180 $X=616900 $Y=633100
X100 2312 2 1 2405 BUF1 $T=618140 557880 1 0 $X=618140 $Y=552460
X101 2293 2 1 2413 BUF1 $T=618140 648600 1 0 $X=618140 $Y=643180
X102 2364 2 1 2404 BUF1 $T=618760 668760 1 0 $X=618760 $Y=663340
X103 2387 2 1 2422 BUF1 $T=621860 638520 1 0 $X=621860 $Y=633100
X104 2379 2 1 2448 BUF1 $T=628060 658680 1 0 $X=628060 $Y=653260
X105 2319 2 1 2444 BUF1 $T=629920 709080 0 0 $X=629920 $Y=708700
X106 2405 2 1 2386 BUF1 $T=630540 567960 0 0 $X=630540 $Y=567580
X107 2402 2 1 2459 BUF1 $T=630540 658680 0 0 $X=630540 $Y=658300
X108 2444 2 1 303 BUF1 $T=633020 709080 0 0 $X=633020 $Y=708700
X109 2405 2 1 2471 BUF1 $T=633640 557880 1 0 $X=633640 $Y=552460
X110 2298 2 1 2461 BUF1 $T=634880 588120 1 0 $X=634880 $Y=582700
X111 2472 2 1 2337 BUF1 $T=637360 608280 0 180 $X=634880 $Y=602860
X112 2387 2 1 2472 BUF1 $T=637360 618360 0 0 $X=637360 $Y=617980
X113 2410 2 1 2494 BUF1 $T=637360 658680 1 0 $X=637360 $Y=653260
X114 2322 2 1 2431 BUF1 $T=637980 567960 1 0 $X=637980 $Y=562540
X115 2422 2 1 2484 BUF1 $T=638600 638520 0 0 $X=638600 $Y=638140
X116 2353 2 1 2492 BUF1 $T=639220 618360 1 0 $X=639220 $Y=612940
X117 2444 2 1 2488 BUF1 $T=639220 699000 1 0 $X=639220 $Y=693580
X118 2461 2 1 300 BUF1 $T=642940 567960 0 180 $X=640460 $Y=562540
X119 2472 2 1 2509 BUF1 $T=649140 618360 1 0 $X=649140 $Y=612940
X120 2444 2 1 2520 BUF1 $T=652860 699000 1 0 $X=652860 $Y=693580
X121 329 2 1 2505 BUF1 $T=654720 709080 0 0 $X=654720 $Y=708700
X122 2461 2 1 2515 BUF1 $T=659060 588120 1 180 $X=656580 $Y=587740
X123 2515 2 1 2584 BUF1 $T=660920 588120 0 0 $X=660920 $Y=587740
X124 329 2 1 2546 BUF1 $T=661540 709080 0 0 $X=661540 $Y=708700
X125 2520 2 1 342 BUF1 $T=670220 709080 1 0 $X=670220 $Y=703660
X126 2520 2 1 2580 BUF1 $T=671460 699000 0 0 $X=671460 $Y=698620
X127 2618 2 1 2621 BUF1 $T=677660 648600 1 0 $X=677660 $Y=643180
X128 2613 2 1 335 BUF1 $T=682620 567960 0 180 $X=680140 $Y=562540
X129 2627 2 1 2651 BUF1 $T=685720 608280 1 0 $X=685720 $Y=602860
X130 2657 2 1 2736 BUF1 $T=699980 567960 0 0 $X=699980 $Y=567580
X131 2656 2 1 2765 BUF1 $T=708040 618360 1 0 $X=708040 $Y=612940
X132 379 2 1 2800 BUF1 $T=719820 709080 0 0 $X=719820 $Y=708700
X133 366 2 1 2900 BUF1 $T=721680 709080 1 0 $X=721680 $Y=703660
X134 2915 2 1 2921 BUF1 $T=725400 709080 0 0 $X=725400 $Y=708700
X135 2925 2 1 2943 BUF1 $T=729120 588120 0 0 $X=729120 $Y=587740
X136 2949 2 1 405 BUF1 $T=732840 719160 1 0 $X=732840 $Y=713740
X137 2673 2 1 3005 BUF1 $T=737180 588120 0 0 $X=737180 $Y=587740
X138 2837 2 1 2987 BUF1 $T=737180 608280 1 0 $X=737180 $Y=602860
X139 2673 2 1 2986 BUF1 $T=738420 588120 1 0 $X=738420 $Y=582700
X140 2949 2 1 3014 BUF1 $T=738420 699000 1 0 $X=738420 $Y=693580
X141 2736 2 1 3045 BUF1 $T=740900 567960 0 0 $X=740900 $Y=567580
X142 367 2 1 3068 BUF1 $T=746480 719160 1 0 $X=746480 $Y=713740
X143 2741 2 1 427 BUF1 $T=759500 699000 1 0 $X=759500 $Y=693580
X144 2671 2 1 3191 BUF1 $T=766320 588120 1 0 $X=766320 $Y=582700
X145 456 2 1 3544 BUF1 $T=820260 699000 1 0 $X=820260 $Y=693580
X146 3547 2 1 3562 BUF1 $T=827080 638520 1 0 $X=827080 $Y=633100
X147 3690 2 1 3700 BUF1 $T=858700 668760 1 0 $X=858700 $Y=663340
X148 3718 2 1 3690 BUF1 $T=864280 668760 1 0 $X=864280 $Y=663340
X149 3830 2 1 3862 BUF1 $T=890320 688920 0 0 $X=890320 $Y=688540
X150 3926 2 1 3929 BUF1 $T=897140 567960 1 0 $X=897140 $Y=562540
X151 589 2 1 4182 BUF1 $T=940540 557880 1 0 $X=940540 $Y=552460
X152 4185 2 1 4047 BUF1 $T=942400 658680 0 0 $X=942400 $Y=658300
X153 3718 2 1 3711 BUF1 $T=947360 638520 1 0 $X=947360 $Y=633100
X154 4185 2 1 4239 BUF1 $T=957900 658680 1 0 $X=957900 $Y=653260
X155 4255 2 1 4202 BUF1 $T=962240 557880 1 180 $X=959760 $Y=557500
X156 4205 2 1 4252 BUF1 $T=968440 578040 0 180 $X=965960 $Y=572620
X157 4295 2 1 4273 BUF1 $T=972160 588120 1 180 $X=969680 $Y=587740
X158 4239 2 1 4313 BUF1 $T=982080 638520 1 0 $X=982080 $Y=633100
X159 4252 2 1 4295 BUF1 $T=984560 578040 1 0 $X=984560 $Y=572620
X160 4295 2 1 4343 BUF1 $T=985180 588120 1 0 $X=985180 $Y=582700
X161 4330 2 1 4359 BUF1 $T=995100 547800 1 0 $X=995100 $Y=542380
X162 641 2 1 4407 BUF1 $T=1015560 709080 0 0 $X=1015560 $Y=708700
X163 4406 2 1 4387 BUF1 $T=1023000 678840 1 180 $X=1020520 $Y=678460
X164 638 2 1 4428 BUF1 $T=1021760 578040 0 0 $X=1021760 $Y=577660
X165 4406 2 1 4449 BUF1 $T=1025480 678840 0 0 $X=1025480 $Y=678460
X166 4452 2 1 4406 BUF1 $T=1029820 688920 0 180 $X=1027340 $Y=683500
X167 4437 2 1 4455 BUF1 $T=1032920 628440 1 180 $X=1030440 $Y=628060
X168 4427 2 1 4409 BUF1 $T=1034160 578040 0 180 $X=1031680 $Y=572620
X169 4455 2 1 4410 BUF1 $T=1037880 618360 0 180 $X=1035400 $Y=612940
X170 638 2 1 648 BUF1 $T=1037260 567960 1 0 $X=1037260 $Y=562540
X171 4508 2 1 4478 BUF1 $T=1058340 648600 1 180 $X=1055860 $Y=648220
X172 4487 2 1 4517 BUF1 $T=1056480 688920 1 0 $X=1056480 $Y=683500
X173 4475 2 1 4509 BUF1 $T=1065780 699000 1 180 $X=1063300 $Y=698620
X174 4523 2 1 655 BUF1 $T=1065160 547800 1 0 $X=1065160 $Y=542380
X175 4508 2 1 4541 BUF1 $T=1065780 648600 0 0 $X=1065780 $Y=648220
X176 4541 2 1 4536 BUF1 $T=1070740 648600 0 0 $X=1070740 $Y=648220
X177 4523 2 1 656 BUF1 $T=1076320 557880 1 0 $X=1076320 $Y=552460
X178 4569 2 1 4568 BUF1 $T=1089960 578040 1 0 $X=1089960 $Y=572620
X179 4618 2 1 4597 BUF1 $T=1111660 608280 0 180 $X=1109180 $Y=602860
X180 858 3 834 2 1 917 QDFFRBN $T=301940 567960 0 0 $X=301940 $Y=567580
X181 924 3 834 2 1 1009 QDFFRBN $T=314340 567960 0 0 $X=314340 $Y=567580
X182 33 11 942 2 1 953 QDFFRBN $T=333560 699000 1 180 $X=321780 $Y=698620
X183 1014 3 985 2 1 1096 QDFFRBN $T=332320 567960 0 0 $X=332320 $Y=567580
X184 1068 11 942 2 1 1043 QDFFRBN $T=347200 688920 1 180 $X=335420 $Y=688540
X185 1056 3 985 2 1 1123 QDFFRBN $T=337280 578040 1 0 $X=337280 $Y=572620
X186 1140 11 1083 2 1 1110 QDFFRBN $T=360840 688920 0 180 $X=349060 $Y=683500
X187 1168 3 985 2 1 1192 QDFFRBN $T=374480 578040 0 180 $X=362700 $Y=572620
X188 1198 11 1083 2 1 1196 QDFFRBN $T=374480 688920 0 180 $X=362700 $Y=683500
X189 1338 11 1303 2 1 977 QDFFRBN $T=388740 668760 1 180 $X=376960 $Y=668380
X190 1286 11 1303 2 1 1333 QDFFRBN $T=376960 678840 0 0 $X=376960 $Y=678460
X191 1343 11 1303 2 1 914 QDFFRBN $T=389360 678840 0 180 $X=377580 $Y=673420
X192 1238 3 1358 2 1 1370 QDFFRBN $T=382540 567960 0 0 $X=382540 $Y=567580
X193 1346 3 1358 2 1 1392 QDFFRBN $T=388120 567960 1 0 $X=388120 $Y=562540
X194 1407 11 1303 2 1 963 QDFFRBN $T=401760 668760 1 180 $X=389980 $Y=668380
X195 1411 11 1303 2 1 932 QDFFRBN $T=402380 678840 0 180 $X=390600 $Y=673420
X196 1451 3 1358 2 1 1383 QDFFRBN $T=409200 557880 1 180 $X=397420 $Y=557500
X197 1402 3 1434 2 1 1455 QDFFRBN $T=398660 578040 1 0 $X=398660 $Y=572620
X198 1454 11 1422 2 1 1001 QDFFRBN $T=411680 658680 1 180 $X=399900 $Y=658300
X199 1457 3 1415 2 1 1313 QDFFRBN $T=413540 598200 0 180 $X=401760 $Y=592780
X200 1449 11 1303 2 1 1401 QDFFRBN $T=413540 668760 1 180 $X=401760 $Y=668380
X201 1456 3 1434 2 1 1425 QDFFRBN $T=416020 567960 1 180 $X=404240 $Y=567580
X202 1498 3 1358 2 1 1457 QDFFRBN $T=422840 557880 1 180 $X=411060 $Y=557500
X203 1512 3 1481 2 1 1462 QDFFRBN $T=424080 588120 1 180 $X=412300 $Y=587740
X204 1470 3 1434 2 1 1529 QDFFRBN $T=412920 578040 1 0 $X=412920 $Y=572620
X205 1462 11 1422 2 1 1468 QDFFRBN $T=424700 658680 1 180 $X=412920 $Y=658300
X206 1482 3 103 2 1 1533 QDFFRBN $T=415400 547800 1 0 $X=415400 $Y=542380
X207 1485 3 1481 2 1 1491 QDFFRBN $T=418500 588120 1 0 $X=418500 $Y=582700
X208 1413 3 103 2 1 1551 QDFFRBN $T=419120 567960 1 0 $X=419120 $Y=562540
X209 1528 3 1549 2 1 1586 QDFFRBN $T=424700 557880 0 0 $X=424700 $Y=557500
X210 1575 11 1422 2 1 104 QDFFRBN $T=436480 658680 1 180 $X=424700 $Y=658300
X211 1537 3 1549 2 1 1575 QDFFRBN $T=427180 578040 1 0 $X=427180 $Y=572620
X212 1609 116 103 2 1 109 QDFFRBN $T=440200 547800 0 180 $X=428420 $Y=542380
X213 1606 11 1568 2 1 1523 QDFFRBN $T=442060 658680 0 180 $X=430280 $Y=653260
X214 1592 116 1481 2 1 1472 QDFFRBN $T=442680 588120 0 180 $X=430900 $Y=582700
X215 1546 11 1568 2 1 1616 QDFFRBN $T=430900 648600 0 0 $X=430900 $Y=648220
X216 1594 116 1549 2 1 1554 QDFFRBN $T=443300 578040 1 180 $X=431520 $Y=577660
X217 1628 11 1568 2 1 1131 QDFFRBN $T=446400 648600 0 180 $X=434620 $Y=643180
X218 1621 116 1358 2 1 1592 QDFFRBN $T=450120 557880 1 180 $X=438340 $Y=557500
X219 1644 116 1358 2 1 1597 QDFFRBN $T=450740 567960 0 180 $X=438960 $Y=562540
X220 1619 116 1641 2 1 1673 QDFFRBN $T=442680 598200 1 0 $X=442680 $Y=592780
X221 1624 116 1641 2 1 1606 QDFFRBN $T=443920 578040 0 0 $X=443920 $Y=577660
X222 1665 11 1568 2 1 1471 QDFFRBN $T=455700 648600 1 180 $X=443920 $Y=648220
X223 1674 11 1635 2 1 989 QDFFRBN $T=455700 668760 0 180 $X=443920 $Y=663340
X224 1668 11 1635 2 1 974 QDFFRBN $T=456320 658680 1 180 $X=444540 $Y=658300
X225 1643 116 1679 2 1 1693 QDFFRBN $T=448880 547800 1 0 $X=448880 $Y=542380
X226 1645 116 1679 2 1 1689 QDFFRBN $T=448880 567960 0 0 $X=448880 $Y=567580
X227 1633 11 1680 2 1 1692 QDFFRBN $T=448880 608280 1 0 $X=448880 $Y=602860
X228 1591 116 1641 2 1 1696 QDFFRBN $T=449500 588120 1 0 $X=449500 $Y=582700
X229 1652 11 1680 2 1 1714 QDFFRBN $T=450740 608280 0 0 $X=450740 $Y=607900
X230 1654 11 1680 2 1 1698 QDFFRBN $T=451360 618360 1 0 $X=451360 $Y=612940
X231 1739 11 1680 2 1 1109 QDFFRBN $T=468100 628440 1 180 $X=456320 $Y=628060
X232 1634 11 1635 2 1 1732 QDFFRBN $T=456320 658680 1 0 $X=456320 $Y=653260
X233 1687 11 1635 2 1 1672 QDFFRBN $T=468100 668760 0 180 $X=456320 $Y=663340
X234 1726 11 1691 2 1 1677 QDFFRBN $T=468100 678840 1 180 $X=456320 $Y=678460
X235 1663 11 1676 2 1 1724 QDFFRBN $T=456940 648600 0 0 $X=456940 $Y=648220
X236 1682 11 1691 2 1 1722 QDFFRBN $T=456940 678840 1 0 $X=456940 $Y=673420
X237 1578 11 1720 2 1 1729 QDFFRBN $T=457560 628440 1 0 $X=457560 $Y=623020
X238 1681 11 1680 2 1 1725 QDFFRBN $T=459420 618360 0 0 $X=459420 $Y=617980
X239 1752 116 143 2 1 138 QDFFRBN $T=474300 547800 0 180 $X=462520 $Y=542380
X240 140 11 1757 2 1 1776 QDFFRBN $T=463760 699000 1 0 $X=463760 $Y=693580
X241 1716 11 1764 2 1 1727 QDFFRBN $T=464380 688920 0 0 $X=464380 $Y=688540
X242 1811 1791 1676 2 1 1741 QDFFRBN $T=480500 658680 1 180 $X=468720 $Y=658300
X243 1802 1791 1691 2 1 1745 QDFFRBN $T=481120 668760 0 180 $X=469340 $Y=663340
X244 1804 152 1691 2 1 1750 QDFFRBN $T=481740 678840 0 180 $X=469960 $Y=673420
X245 1805 152 1691 2 1 1742 QDFFRBN $T=481740 678840 1 180 $X=469960 $Y=678460
X246 1808 1791 1720 2 1 1536 QDFFRBN $T=482360 628440 0 180 $X=470580 $Y=623020
X247 1809 1791 1720 2 1 1339 QDFFRBN $T=482360 628440 1 180 $X=470580 $Y=628060
X248 1810 1791 1720 2 1 1752 QDFFRBN $T=482360 638520 0 180 $X=470580 $Y=633100
X249 1801 1791 1676 2 1 1665 QDFFRBN $T=482360 648600 1 180 $X=470580 $Y=648220
X250 1816 1791 1720 2 1 1189 QDFFRBN $T=482980 638520 1 180 $X=471200 $Y=638140
X251 1761 11 1757 2 1 1828 QDFFRBN $T=471820 709080 1 0 $X=471820 $Y=703660
X252 1846 11 1757 2 1 1779 QDFFRBN $T=487320 699000 0 180 $X=475540 $Y=693580
X253 1803 152 1764 2 1 1859 QDFFRBN $T=479260 688920 1 0 $X=479260 $Y=683500
X254 1821 1791 1842 2 1 1873 QDFFRBN $T=481740 618360 0 0 $X=481740 $Y=617980
X255 1872 1791 1842 2 1 1824 QDFFRBN $T=494140 638520 0 180 $X=482360 $Y=633100
X256 1866 1791 1676 2 1 1825 QDFFRBN $T=494140 658680 1 180 $X=482360 $Y=658300
X257 1827 1791 1842 2 1 1874 QDFFRBN $T=482980 628440 1 0 $X=482980 $Y=623020
X258 1832 1791 1842 2 1 1881 QDFFRBN $T=483600 598200 0 0 $X=483600 $Y=597820
X259 1834 11 151 2 1 169 QDFFRBN $T=483600 719160 1 0 $X=483600 $Y=713740
X260 1837 116 1679 2 1 1887 QDFFRBN $T=484840 578040 0 0 $X=484840 $Y=577660
X261 1904 1791 1842 2 1 1836 QDFFRBN $T=496620 618360 0 180 $X=484840 $Y=612940
X262 1844 116 1679 2 1 1870 QDFFRBN $T=485460 567960 1 0 $X=485460 $Y=562540
X263 1813 116 1679 2 1 1892 QDFFRBN $T=486080 557880 0 0 $X=486080 $Y=557500
X264 1897 1791 1851 2 1 1855 QDFFRBN $T=500340 658680 0 180 $X=488560 $Y=653260
X265 1867 152 175 2 1 1914 QDFFRBN $T=491660 709080 1 0 $X=491660 $Y=703660
X266 1871 116 1896 2 1 1900 QDFFRBN $T=492280 578040 1 0 $X=492280 $Y=572620
X267 1912 152 1764 2 1 1869 QDFFRBN $T=504060 688920 0 180 $X=492280 $Y=683500
X268 1923 116 1896 2 1 1885 QDFFRBN $T=507160 598200 1 180 $X=495380 $Y=597820
X269 1899 152 151 2 1 171 QDFFRBN $T=507160 719160 0 180 $X=495380 $Y=713740
X270 1929 1791 1863 2 1 1886 QDFFRBN $T=507780 628440 1 180 $X=496000 $Y=628060
X271 1919 1791 1851 2 1 1890 QDFFRBN $T=509640 658680 1 180 $X=497860 $Y=658300
X272 1905 152 175 2 1 1948 QDFFRBN $T=500340 699000 0 0 $X=500340 $Y=698620
X273 1925 1791 1851 2 1 1907 QDFFRBN $T=512740 668760 0 180 $X=500960 $Y=663340
X274 1909 116 1896 2 1 1944 QDFFRBN $T=501580 578040 0 0 $X=501580 $Y=577660
X275 1957 152 175 2 1 1913 QDFFRBN $T=514600 709080 1 180 $X=502820 $Y=708700
X276 1916 1791 1863 2 1 1962 QDFFRBN $T=503440 608280 0 0 $X=503440 $Y=607900
X277 1917 1791 1863 2 1 1956 QDFFRBN $T=503440 618360 0 0 $X=503440 $Y=617980
X278 1921 116 1952 2 1 1941 QDFFRBN $T=504680 578040 1 0 $X=504680 $Y=572620
X279 1936 152 1764 2 1 1920 QDFFRBN $T=517080 688920 0 180 $X=505300 $Y=683500
X280 1965 1791 1851 2 1 1924 QDFFRBN $T=517700 658680 0 180 $X=505920 $Y=653260
X281 1933 116 165 2 1 1976 QDFFRBN $T=507780 547800 0 0 $X=507780 $Y=547420
X282 1981 1791 1863 2 1 1932 QDFFRBN $T=519560 628440 1 180 $X=507780 $Y=628060
X283 1947 152 1986 2 1 2006 QDFFRBN $T=510880 699000 1 0 $X=510880 $Y=693580
X284 1951 116 1952 2 1 1977 QDFFRBN $T=511500 567960 0 0 $X=511500 $Y=567580
X285 1964 1791 2002 2 1 1993 QDFFRBN $T=514600 628440 1 0 $X=514600 $Y=623020
X286 1969 152 2007 2 1 2017 QDFFRBN $T=515220 709080 0 0 $X=515220 $Y=708700
X287 1999 116 1952 2 1 1970 QDFFRBN $T=527620 578040 1 180 $X=515840 $Y=577660
X288 1973 1791 2009 2 1 2014 QDFFRBN $T=515840 668760 1 0 $X=515840 $Y=663340
X289 1980 116 1952 2 1 2025 QDFFRBN $T=517700 567960 1 0 $X=517700 $Y=562540
X290 1967 152 1986 2 1 2029 QDFFRBN $T=517700 678840 0 0 $X=517700 $Y=678460
X291 1975 1791 1851 2 1 2016 QDFFRBN $T=518320 658680 1 0 $X=518320 $Y=653260
X292 1991 116 1896 2 1 2044 QDFFRBN $T=520180 598200 0 0 $X=520180 $Y=597820
X293 2030 152 1986 2 1 1995 QDFFRBN $T=533200 678840 0 180 $X=521420 $Y=673420
X294 2001 152 1986 2 1 2022 QDFFRBN $T=523280 688920 1 0 $X=523280 $Y=683500
X295 2045 152 2007 2 1 1983 QDFFRBN $T=535060 709080 0 180 $X=523280 $Y=703660
X296 2015 1791 2002 2 1 2012 QDFFRBN $T=537540 618360 1 180 $X=525760 $Y=617980
X297 2023 1791 2002 2 1 2047 QDFFRBN $T=527000 628440 0 0 $X=527000 $Y=628060
X298 2005 1791 2052 2 1 2072 QDFFRBN $T=527000 648600 0 0 $X=527000 $Y=648220
X299 2027 116 2055 2 1 2042 QDFFRBN $T=527620 608280 1 0 $X=527620 $Y=602860
X300 2040 1791 2002 2 1 2018 QDFFRBN $T=539400 628440 0 180 $X=527620 $Y=623020
X301 2065 152 2007 2 1 2026 QDFFRBN $T=539400 709080 1 180 $X=527620 $Y=708700
X302 2066 116 196 2 1 2031 QDFFRBN $T=541880 547800 0 180 $X=530100 $Y=542380
X303 2078 116 2046 2 1 2035 QDFFRBN $T=542500 567960 0 180 $X=530720 $Y=562540
X304 2037 1791 2067 2 1 2059 QDFFRBN $T=530720 638520 0 0 $X=530720 $Y=638140
X305 2038 152 2009 2 1 2083 QDFFRBN $T=530720 678840 0 0 $X=530720 $Y=678460
X306 2098 1791 2067 2 1 2056 QDFFRBN $T=547460 638520 0 180 $X=535680 $Y=633100
X307 2054 1791 2088 2 1 2060 QDFFRBN $T=538780 618360 1 0 $X=538780 $Y=612940
X308 2071 1791 2088 2 1 2099 QDFFRBN $T=538780 618360 0 0 $X=538780 $Y=617980
X309 2070 116 2046 2 1 2112 QDFFRBN $T=539400 578040 1 0 $X=539400 $Y=572620
X310 2109 1791 2055 2 1 2076 QDFFRBN $T=552420 608280 0 180 $X=540640 $Y=602860
X311 2097 152 2009 2 1 2086 QDFFRBN $T=554280 678840 1 180 $X=542500 $Y=678460
X312 2092 1791 2052 2 1 2126 QDFFRBN $T=543120 658680 0 0 $X=543120 $Y=658300
X313 2075 152 243 2 1 2127 QDFFRBN $T=544360 719160 1 0 $X=544360 $Y=713740
X314 2089 152 2108 2 1 2122 QDFFRBN $T=544980 699000 0 0 $X=544980 $Y=698620
X315 2101 152 243 2 1 2091 QDFFRBN $T=556760 709080 1 180 $X=544980 $Y=708700
X316 2100 1791 2067 2 1 2140 QDFFRBN $T=546840 648600 1 0 $X=546840 $Y=643180
X317 2135 250 2046 2 1 2102 QDFFRBN $T=559240 567960 0 180 $X=547460 $Y=562540
X318 2139 1791 2067 2 1 2104 QDFFRBN $T=559860 628440 0 180 $X=548080 $Y=623020
X319 2106 1791 2067 2 1 2143 QDFFRBN $T=548080 638520 1 0 $X=548080 $Y=633100
X320 2137 152 2108 2 1 2105 QDFFRBN $T=559860 688920 0 180 $X=548080 $Y=683500
X321 2136 1791 2055 2 1 2107 QDFFRBN $T=560480 598200 1 180 $X=548700 $Y=597820
X322 2155 250 2046 2 1 2114 QDFFRBN $T=562340 567960 1 180 $X=550560 $Y=567580
X323 2113 152 2146 2 1 2115 QDFFRBN $T=551180 678840 1 0 $X=551180 $Y=673420
X324 2168 250 2123 2 1 2118 QDFFRBN $T=563580 588120 0 180 $X=551800 $Y=582700
X325 2119 1791 2148 2 1 2162 QDFFRBN $T=551800 618360 1 0 $X=551800 $Y=612940
X326 2134 1791 2146 2 1 2182 QDFFRBN $T=556760 658680 0 0 $X=556760 $Y=658300
X327 2138 152 255 2 1 2196 QDFFRBN $T=559240 709080 0 0 $X=559240 $Y=708700
X328 2152 152 2108 2 1 2195 QDFFRBN $T=559860 688920 1 0 $X=559860 $Y=683500
X329 2156 1791 2186 2 1 2178 QDFFRBN $T=560480 648600 1 0 $X=560480 $Y=643180
X330 2157 1791 2186 2 1 2184 QDFFRBN $T=561100 638520 1 0 $X=561100 $Y=633100
X331 2161 1791 2148 2 1 2202 QDFFRBN $T=561720 628440 1 0 $X=561720 $Y=623020
X332 2190 1791 2172 2 1 2163 QDFFRBN $T=574740 678840 0 180 $X=562960 $Y=673420
X333 2144 152 255 2 1 2200 QDFFRBN $T=562960 699000 0 0 $X=562960 $Y=698620
X334 256 152 255 2 1 2210 QDFFRBN $T=563580 719160 1 0 $X=563580 $Y=713740
X335 2213 250 260 2 1 2169 QDFFRBN $T=576600 567960 0 180 $X=564820 $Y=562540
X336 1815 1791 2148 2 1 2223 QDFFRBN $T=565440 618360 1 0 $X=565440 $Y=612940
X337 2183 1791 2146 2 1 2221 QDFFRBN $T=566680 668760 0 0 $X=566680 $Y=668380
X338 2216 1791 2164 2 1 2185 QDFFRBN $T=580320 598200 0 180 $X=568540 $Y=592780
X339 2222 1791 2123 2 1 2192 QDFFRBN $T=581560 588120 1 180 $X=569780 $Y=587740
X340 2231 1791 2186 2 1 2193 QDFFRBN $T=581560 628440 1 180 $X=569780 $Y=628060
X341 266 1791 2186 2 1 259 QDFFRBN $T=581560 638520 1 180 $X=569780 $Y=638140
X342 2189 1791 2146 2 1 2198 QDFFRBN $T=570400 658680 0 0 $X=570400 $Y=658300
X343 2199 152 2172 2 1 2239 QDFFRBN $T=572260 688920 1 0 $X=572260 $Y=683500
X344 2240 271 2146 2 1 2206 QDFFRBN $T=585280 668760 0 180 $X=573500 $Y=663340
X345 2243 250 260 2 1 2204 QDFFRBN $T=585900 557880 0 180 $X=574120 $Y=552460
X346 1807 1791 2237 2 1 2254 QDFFRBN $T=574120 598200 0 0 $X=574120 $Y=597820
X347 2208 152 2226 2 1 2251 QDFFRBN $T=574120 699000 1 0 $X=574120 $Y=693580
X348 2215 1791 2148 2 1 2259 QDFFRBN $T=575980 618360 0 0 $X=575980 $Y=617980
X349 265 152 261 2 1 2257 QDFFRBN $T=576600 719160 1 0 $X=576600 $Y=713740
X350 2225 250 2233 2 1 2272 QDFFRBN $T=578460 567960 1 0 $X=578460 $Y=562540
X351 2244 250 2233 2 1 2217 QDFFRBN $T=590240 578040 1 180 $X=578460 $Y=577660
X352 2269 271 2207 2 1 2230 QDFFRBN $T=591480 648600 0 180 $X=579700 $Y=643180
X353 2232 152 2261 2 1 2279 QDFFRBN $T=580320 678840 1 0 $X=580320 $Y=673420
X354 2245 152 2261 2 1 2297 QDFFRBN $T=584660 678840 0 0 $X=584660 $Y=678460
X355 2294 2290 2237 2 1 2246 QDFFRBN $T=597060 608280 0 180 $X=585280 $Y=602860
X356 1857 250 2233 2 1 2307 QDFFRBN $T=586520 578040 1 0 $X=586520 $Y=572620
X357 2265 271 2293 2 1 2318 QDFFRBN $T=588380 658680 0 0 $X=588380 $Y=658300
X358 2302 271 2226 2 1 2264 QDFFRBN $T=600780 699000 0 180 $X=589000 $Y=693580
X359 1848 250 2233 2 1 2323 QDFFRBN $T=589620 588120 1 0 $X=589620 $Y=582700
X360 2263 271 277 2 1 2324 QDFFRBN $T=589620 709080 0 0 $X=589620 $Y=708700
X361 2314 250 2233 2 1 2270 QDFFRBN $T=602020 567960 1 180 $X=590240 $Y=567580
X362 2274 250 273 2 1 2326 QDFFRBN $T=590860 547800 1 0 $X=590860 $Y=542380
X363 2275 250 280 2 1 2327 QDFFRBN $T=590860 557880 0 0 $X=590860 $Y=557500
X364 2287 2290 2237 2 1 2321 QDFFRBN $T=592720 608280 0 0 $X=592720 $Y=607900
X365 2329 2290 2266 2 1 2285 QDFFRBN $T=604500 638520 0 180 $X=592720 $Y=633100
X366 2289 250 2320 2 1 2283 QDFFRBN $T=593340 578040 0 0 $X=593340 $Y=577660
X367 2292 271 2293 2 1 2336 QDFFRBN $T=593340 668760 1 0 $X=593340 $Y=663340
X368 2301 271 2261 2 1 2352 QDFFRBN $T=596440 688920 0 0 $X=596440 $Y=688540
X369 2348 271 2316 2 1 2304 QDFFRBN $T=609460 668760 1 180 $X=597680 $Y=668380
X370 2308 271 2261 2 1 2346 QDFFRBN $T=598300 688920 1 0 $X=598300 $Y=683500
X371 2313 250 2320 2 1 2363 QDFFRBN $T=599540 578040 1 0 $X=599540 $Y=572620
X372 2347 2290 2266 2 1 2317 QDFFRBN $T=613800 638520 1 180 $X=602020 $Y=638140
X373 2367 2290 2316 2 1 2325 QDFFRBN $T=614420 658680 1 180 $X=602640 $Y=658300
X374 2333 271 277 2 1 2371 QDFFRBN $T=603260 709080 0 0 $X=603260 $Y=708700
X375 286 250 280 2 1 2381 QDFFRBN $T=603880 547800 1 0 $X=603880 $Y=542380
X376 2335 250 280 2 1 2368 QDFFRBN $T=603880 557880 0 0 $X=603880 $Y=557500
X377 1830 250 2360 2 1 2377 QDFFRBN $T=603880 567960 0 0 $X=603880 $Y=567580
X378 2310 271 277 2 1 293 QDFFRBN $T=603880 719160 1 0 $X=603880 $Y=713740
X379 2339 2290 2353 2 1 2362 QDFFRBN $T=605120 608280 0 0 $X=605120 $Y=607900
X380 2374 2290 2353 2 1 2341 QDFFRBN $T=617520 628440 1 180 $X=605740 $Y=628060
X381 2343 250 280 2 1 2389 QDFFRBN $T=606360 557880 1 0 $X=606360 $Y=552460
X382 2393 2290 2320 2 1 2344 QDFFRBN $T=619380 578040 1 180 $X=607600 $Y=577660
X383 2380 271 2316 2 1 2358 QDFFRBN $T=621240 668760 1 180 $X=609460 $Y=668380
X384 2359 271 296 2 1 2420 QDFFRBN $T=611940 699000 1 0 $X=611940 $Y=693580
X385 2365 271 296 2 1 2417 QDFFRBN $T=611940 709080 1 0 $X=611940 $Y=703660
X386 2397 2290 2353 2 1 2366 QDFFRBN $T=626200 618360 0 180 $X=614420 $Y=612940
X387 2383 2290 2413 2 1 2429 QDFFRBN $T=615660 638520 0 0 $X=615660 $Y=638140
X388 2426 271 2316 2 1 2382 QDFFRBN $T=627440 678840 0 180 $X=615660 $Y=673420
X389 2385 250 300 2 1 2433 QDFFRBN $T=616280 557880 0 0 $X=616280 $Y=557500
X390 2388 271 296 2 1 2439 QDFFRBN $T=616280 709080 0 0 $X=616280 $Y=708700
X391 2395 2290 2360 2 1 2441 QDFFRBN $T=617520 608280 0 0 $X=617520 $Y=607900
X392 2398 2290 2353 2 1 2428 QDFFRBN $T=618760 628440 0 0 $X=618760 $Y=628060
X393 2414 271 2293 2 1 2463 QDFFRBN $T=621860 668760 1 0 $X=621860 $Y=663340
X394 2460 2290 2360 2 1 2416 QDFFRBN $T=634260 598200 0 180 $X=622480 $Y=592780
X395 2401 271 2316 2 1 2442 QDFFRBN $T=622480 668760 0 0 $X=622480 $Y=668380
X396 2419 2290 2293 2 1 2466 QDFFRBN $T=623100 648600 1 0 $X=623100 $Y=643180
X397 2457 271 296 2 1 2423 QDFFRBN $T=636120 709080 0 180 $X=624340 $Y=703660
X398 2453 271 296 2 1 2425 QDFFRBN $T=636740 699000 0 180 $X=624960 $Y=693580
X399 2467 2290 2353 2 1 2436 QDFFRBN $T=639220 618360 0 180 $X=627440 $Y=612940
X400 2445 250 300 2 1 2458 QDFFRBN $T=629300 557880 0 0 $X=629300 $Y=557500
X401 2446 250 2461 2 1 2486 QDFFRBN $T=629300 578040 1 0 $X=629300 $Y=572620
X402 2479 250 300 2 1 2447 QDFFRBN $T=641700 547800 0 180 $X=629920 $Y=542380
X403 2454 2290 2461 2 1 2440 QDFFRBN $T=641700 588120 1 180 $X=629920 $Y=587740
X404 2496 271 2462 2 1 2449 QDFFRBN $T=641700 678840 0 180 $X=629920 $Y=673420
X405 2452 271 2462 2 1 2490 QDFFRBN $T=630540 678840 0 0 $X=630540 $Y=678460
X406 2456 271 2462 2 1 2499 QDFFRBN $T=631780 688920 0 0 $X=631780 $Y=688540
X407 2450 2290 2413 2 1 2465 QDFFRBN $T=646040 638520 0 180 $X=634260 $Y=633100
X408 2470 2290 2492 2 1 2513 QDFFRBN $T=634880 608280 0 0 $X=634880 $Y=607900
X409 2493 2290 2413 2 1 2469 QDFFRBN $T=646660 648600 0 180 $X=634880 $Y=643180
X410 2475 271 2505 2 1 2518 QDFFRBN $T=636740 709080 1 0 $X=636740 $Y=703660
X411 2480 2290 2492 2 1 2521 QDFFRBN $T=638600 628440 1 0 $X=638600 $Y=623020
X412 2481 2290 2461 2 1 2519 QDFFRBN $T=639220 588120 1 0 $X=639220 $Y=582700
X413 2482 2290 2515 2 1 2504 QDFFRBN $T=639220 598200 0 0 $X=639220 $Y=597820
X414 2489 2290 2413 2 1 2536 QDFFRBN $T=641080 638520 0 0 $X=641080 $Y=638140
X415 2491 250 2461 2 1 2553 QDFFRBN $T=641700 578040 1 0 $X=641700 $Y=572620
X416 2495 271 2462 2 1 2531 QDFFRBN $T=641700 668760 0 0 $X=641700 $Y=668380
X417 2497 271 2462 2 1 2545 QDFFRBN $T=641700 678840 1 0 $X=641700 $Y=673420
X418 2524 250 321 2 1 317 QDFFRBN $T=655340 547800 0 180 $X=643560 $Y=542380
X419 2528 2290 2515 2 1 2506 QDFFRBN $T=656580 598200 0 180 $X=644800 $Y=592780
X420 2507 2290 2413 2 1 2517 QDFFRBN $T=644800 648600 0 0 $X=644800 $Y=648220
X421 2500 271 2505 2 1 2562 QDFFRBN $T=645420 699000 0 0 $X=645420 $Y=698620
X422 2512 271 2546 2 1 2533 QDFFRBN $T=646040 688920 0 0 $X=646040 $Y=688540
X423 2514 2290 2413 2 1 2563 QDFFRBN $T=646660 638520 1 0 $X=646660 $Y=633100
X424 2559 2290 2515 2 1 2529 QDFFRBN $T=663400 598200 1 180 $X=651620 $Y=597820
X425 2548 2290 2492 2 1 2523 QDFFRBN $T=664020 608280 1 180 $X=652240 $Y=607900
X426 2537 2290 2492 2 1 2569 QDFFRBN $T=652240 618360 0 0 $X=652240 $Y=617980
X427 2592 271 2505 2 1 2532 QDFFRBN $T=665880 709080 0 180 $X=654100 $Y=703660
X428 2547 250 335 2 1 332 QDFFRBN $T=656580 547800 0 0 $X=656580 $Y=547420
X429 2544 2290 2584 2 1 2554 QDFFRBN $T=656580 588120 1 0 $X=656580 $Y=582700
X430 2558 2290 2584 2 1 2571 QDFFRBN $T=657200 578040 0 0 $X=657200 $Y=577660
X431 2561 271 2546 2 1 2593 QDFFRBN $T=657200 699000 1 0 $X=657200 $Y=693580
X432 2527 250 2584 2 1 2594 QDFFRBN $T=657820 567960 0 0 $X=657820 $Y=567580
X433 2552 271 2557 2 1 2576 QDFFRBN $T=657820 668760 1 0 $X=657820 $Y=663340
X434 2567 250 335 2 1 336 QDFFRBN $T=658440 557880 1 0 $X=658440 $Y=552460
X435 2571 2290 2515 2 1 2615 QDFFRBN $T=658440 598200 1 0 $X=658440 $Y=592780
X436 2541 250 335 2 1 2566 QDFFRBN $T=659060 567960 1 0 $X=659060 $Y=562540
X437 2574 2290 2589 2 1 2598 QDFFRBN $T=659680 618360 1 0 $X=659680 $Y=612940
X438 339 271 329 2 1 2573 QDFFRBN $T=671460 719160 0 180 $X=659680 $Y=713740
X439 2578 250 341 2 1 343 QDFFRBN $T=662780 547800 1 0 $X=662780 $Y=542380
X440 2585 271 2546 2 1 2609 QDFFRBN $T=664020 688920 1 0 $X=664020 $Y=683500
X441 2586 271 2546 2 1 2612 QDFFRBN $T=664020 709080 0 0 $X=664020 $Y=708700
X442 2590 250 2613 2 1 2599 QDFFRBN $T=667740 588120 0 0 $X=667740 $Y=587740
X443 2587 2290 2600 2 1 2603 QDFFRBN $T=667740 658680 0 0 $X=667740 $Y=658300
X444 2591 2290 2557 2 1 2620 QDFFRBN $T=667740 668760 0 0 $X=667740 $Y=668380
X445 2582 2290 2589 2 1 2624 QDFFRBN $T=668360 618360 0 0 $X=668360 $Y=617980
X446 2553 2290 2589 2 1 2639 QDFFRBN $T=671460 608280 0 0 $X=671460 $Y=607900
X447 2468 2290 2621 2 1 2636 QDFFRBN $T=671460 628440 0 0 $X=671460 $Y=628060
X448 2601 250 335 2 1 353 QDFFRBN $T=672080 557880 1 0 $X=672080 $Y=552460
X449 2625 250 341 2 1 344 QDFFRBN $T=686960 547800 0 180 $X=675180 $Y=542380
X450 2607 250 335 2 1 2602 QDFFRBN $T=687580 557880 1 180 $X=675800 $Y=557500
X451 2594 250 2613 2 1 2657 QDFFRBN $T=675800 567960 0 0 $X=675800 $Y=567580
X452 2616 271 2641 2 1 2652 QDFFRBN $T=676420 688920 0 0 $X=676420 $Y=688540
X453 2610 271 357 2 1 360 QDFFRBN $T=677040 719160 1 0 $X=677040 $Y=713740
X454 2623 271 357 2 1 2661 QDFFRBN $T=678900 709080 1 0 $X=678900 $Y=703660
X455 2619 271 2641 2 1 2660 QDFFRBN $T=680760 699000 1 0 $X=680760 $Y=693580
X456 2451 2290 2618 2 1 2662 QDFFRBN $T=681380 648600 1 0 $X=681380 $Y=643180
X457 2418 2290 2618 2 1 2642 QDFFRBN $T=681380 658680 1 0 $X=681380 $Y=653260
X458 2421 2290 2611 2 1 2645 QDFFRBN $T=681380 668760 1 0 $X=681380 $Y=663340
X459 2437 2290 2668 2 1 2697 QDFFRBN $T=685100 628440 0 0 $X=685100 $Y=628060
X460 358 271 2611 2 1 2715 QDFFRBN $T=685720 668760 0 0 $X=685720 $Y=668380
X461 2632 271 2611 2 1 2646 QDFFRBN $T=685720 678840 1 0 $X=685720 $Y=673420
X462 2652 271 2641 2 1 2741 QDFFRBN $T=691300 688920 0 0 $X=691300 $Y=688540
X463 2565 2290 2668 2 1 2727 QDFFRBN $T=694400 638520 1 0 $X=694400 $Y=633100
X464 2392 2290 2668 2 1 2762 QDFFRBN $T=695020 638520 0 0 $X=695020 $Y=638140
X465 2549 2290 2668 2 1 2792 QDFFRBN $T=700600 648600 0 0 $X=700600 $Y=648220
X466 1771 439 443 2 1 446 QDFFRBN $T=791740 547800 1 0 $X=791740 $Y=542380
X467 452 439 457 2 1 3521 QDFFRBN $T=809100 547800 0 0 $X=809100 $Y=547420
X468 1320 439 3538 2 1 3561 QDFFRBN $T=819020 567960 1 0 $X=819020 $Y=562540
X469 1127 439 3538 2 1 3568 QDFFRBN $T=819640 567960 0 0 $X=819640 $Y=567580
X470 1328 439 3538 2 1 3588 QDFFRBN $T=820260 557880 0 0 $X=820260 $Y=557500
X471 1308 439 3538 2 1 3611 QDFFRBN $T=821500 578040 0 0 $X=821500 $Y=577660
X472 3532 465 3562 2 1 3569 QDFFRBN $T=822120 628440 0 0 $X=822120 $Y=628060
X473 462 465 3547 2 1 3575 QDFFRBN $T=822120 648600 1 0 $X=822120 $Y=643180
X474 3534 465 3562 2 1 3581 QDFFRBN $T=823360 638520 0 0 $X=823360 $Y=638140
X475 478 465 3547 2 1 3546 QDFFRBN $T=838860 648600 1 180 $X=827080 $Y=648220
X476 980 439 469 2 1 3615 QDFFRBN $T=828320 547800 0 0 $X=828320 $Y=547420
X477 1304 439 469 2 1 3616 QDFFRBN $T=828940 557880 1 0 $X=828940 $Y=552460
X478 3607 465 3592 2 1 3570 QDFFRBN $T=844440 638520 0 180 $X=832660 $Y=633100
X479 3600 465 3592 2 1 3580 QDFFRBN $T=845680 628440 0 180 $X=833900 $Y=623020
X480 3573 465 3592 2 1 3620 QDFFRBN $T=834520 628440 0 0 $X=834520 $Y=628060
X481 3567 465 3637 2 1 3682 QDFFRBN $T=840100 668760 1 0 $X=840100 $Y=663340
X482 490 465 493 2 1 3709 QDFFRBN $T=848160 719160 1 0 $X=848160 $Y=713740
X483 3683 465 3592 2 1 489 QDFFRBN $T=860560 628440 1 180 $X=848780 $Y=628060
X484 3705 465 493 2 1 3656 QDFFRBN $T=861180 709080 0 180 $X=849400 $Y=703660
X485 3563 465 3690 2 1 3719 QDFFRBN $T=850020 668760 0 0 $X=850020 $Y=668380
X486 3559 465 3700 2 1 3727 QDFFRBN $T=850640 678840 1 0 $X=850640 $Y=673420
X487 3536 465 3690 2 1 3722 QDFFRBN $T=853120 678840 0 0 $X=853120 $Y=678460
X488 3712 465 3592 2 1 492 QDFFRBN $T=866140 628440 0 180 $X=854360 $Y=623020
X489 3689 465 3711 2 1 3725 QDFFRBN $T=854360 699000 1 0 $X=854360 $Y=693580
X490 3717 439 3702 2 1 495 QDFFRBN $T=866760 608280 1 180 $X=854980 $Y=607900
X491 3721 439 3702 2 1 496 QDFFRBN $T=866760 618360 0 180 $X=854980 $Y=612940
X492 3577 465 3690 2 1 3734 QDFFRBN $T=856220 688920 1 0 $X=856220 $Y=683500
X493 3574 465 3711 2 1 3758 QDFFRBN $T=856840 688920 0 0 $X=856840 $Y=688540
X494 3737 439 3702 2 1 494 QDFFRBN $T=869240 608280 0 180 $X=857460 $Y=602860
X495 978 439 3702 2 1 3792 QDFFRBN $T=858080 598200 0 0 $X=858080 $Y=597820
X496 3808 465 3702 2 1 3706 QDFFRBN $T=877300 618360 1 180 $X=865520 $Y=617980
X497 3560 465 3700 2 1 3802 QDFFRBN $T=866140 678840 0 0 $X=866140 $Y=678460
X498 3848 465 3700 2 1 3764 QDFFRBN $T=882880 688920 0 180 $X=871100 $Y=683500
X499 3886 465 3700 2 1 3748 QDFFRBN $T=883500 678840 0 180 $X=871720 $Y=673420
X500 3842 439 3783 2 1 3707 QDFFRBN $T=885980 608280 1 180 $X=874200 $Y=607900
X501 3851 439 3783 2 1 3778 QDFFRBN $T=887220 618360 0 180 $X=875440 $Y=612940
X502 3810 465 3700 2 1 3870 QDFFRBN $T=879160 678840 0 0 $X=879160 $Y=678460
X503 3940 439 3783 2 1 3726 QDFFRBN $T=898380 608280 1 180 $X=886600 $Y=607900
X504 3930 439 3783 2 1 3859 QDFFRBN $T=899620 618360 0 180 $X=887840 $Y=612940
X505 4054 439 3783 2 1 543 QDFFRBN $T=912020 608280 1 180 $X=900240 $Y=607900
X506 4008 439 3783 2 1 544 QDFFRBN $T=912020 618360 0 180 $X=900240 $Y=612940
X507 3996 439 4041 2 1 4048 QDFFRBN $T=908300 608280 1 0 $X=908300 $Y=602860
X508 4073 4080 4041 2 1 3961 QDFFRBN $T=925040 618360 0 180 $X=913260 $Y=612940
X509 4121 4080 4041 2 1 4021 QDFFRBN $T=931860 608280 0 180 $X=920080 $Y=602860
X510 4181 4080 4041 2 1 3986 QDFFRBN $T=943640 608280 0 180 $X=931860 $Y=602860
X511 581 585 4182 2 1 4206 QDFFRBN $T=936200 547800 0 0 $X=936200 $Y=547420
X512 4206 585 589 2 1 583 QDFFRBN $T=948600 547800 0 180 $X=936820 $Y=542380
X513 4208 585 589 2 1 4164 QDFFRBN $T=949220 557880 1 180 $X=937440 $Y=557500
X514 4167 585 4202 2 1 4208 QDFFRBN $T=938060 567960 1 0 $X=938060 $Y=562540
X515 4212 585 4182 2 1 4167 QDFFRBN $T=950460 567960 1 180 $X=938680 $Y=567580
X516 4168 4080 3711 2 1 4198 QDFFRBN $T=939300 598200 1 0 $X=939300 $Y=592780
X517 4063 4080 4205 2 1 4204 QDFFRBN $T=940540 588120 0 0 $X=940540 $Y=587740
X518 4194 4080 4041 2 1 4197 QDFFRBN $T=944260 608280 1 0 $X=944260 $Y=602860
X519 4197 4080 3711 2 1 4235 QDFFRBN $T=944260 608280 0 0 $X=944260 $Y=607900
X520 4198 4080 3711 2 1 4248 QDFFRBN $T=944880 598200 0 0 $X=944880 $Y=597820
X521 4204 4080 4205 2 1 4224 QDFFRBN $T=946120 588120 1 0 $X=946120 $Y=582700
X522 4235 4080 4213 2 1 4203 QDFFRBN $T=957900 618360 0 180 $X=946120 $Y=612940
X523 4203 4080 4213 2 1 4236 QDFFRBN $T=946740 618360 0 0 $X=946740 $Y=617980
X524 4261 585 4202 2 1 4220 QDFFRBN $T=963480 567960 0 180 $X=951700 $Y=562540
X525 4223 585 4252 2 1 4244 QDFFRBN $T=951700 578040 1 0 $X=951700 $Y=572620
X526 4224 585 4202 2 1 4261 QDFFRBN $T=952320 567960 0 0 $X=952320 $Y=567580
X527 4236 4080 4247 2 1 4277 QDFFRBN $T=956040 638520 1 0 $X=956040 $Y=633100
X528 4232 4080 4247 2 1 4292 QDFFRBN $T=956040 638520 0 0 $X=956040 $Y=638140
X529 4244 4080 4273 2 1 4246 QDFFRBN $T=957280 598200 1 0 $X=957280 $Y=592780
X530 4277 4080 4247 2 1 4240 QDFFRBN $T=969060 648600 0 180 $X=957280 $Y=643180
X531 4248 4080 4273 2 1 4284 QDFFRBN $T=957900 598200 0 0 $X=957900 $Y=597820
X532 4240 4080 4247 2 1 4282 QDFFRBN $T=957900 648600 0 0 $X=957900 $Y=648220
X533 4058 585 4205 2 1 4266 QDFFRBN $T=958520 588120 1 0 $X=958520 $Y=582700
X534 3960 585 4205 2 1 4304 QDFFRBN $T=960380 578040 0 0 $X=960380 $Y=577660
X535 4266 585 4255 2 1 4283 QDFFRBN $T=963480 557880 0 0 $X=963480 $Y=557500
X536 4304 585 4255 2 1 4262 QDFFRBN $T=976500 567960 0 180 $X=964720 $Y=562540
X537 4282 4080 4239 2 1 4323 QDFFRBN $T=968440 658680 0 0 $X=968440 $Y=658300
X538 4288 4080 4309 2 1 4281 QDFFRBN $T=969680 628440 1 0 $X=969680 $Y=623020
X539 4292 4080 4313 2 1 4322 QDFFRBN $T=969680 638520 0 0 $X=969680 $Y=638140
X540 4294 585 4252 2 1 4299 QDFFRBN $T=970300 567960 0 0 $X=970300 $Y=567580
X541 4321 4080 4213 2 1 4288 QDFFRBN $T=982080 608280 1 180 $X=970300 $Y=607900
X542 4322 4080 4239 2 1 4291 QDFFRBN $T=982080 648600 0 180 $X=970300 $Y=643180
X543 4316 585 4252 2 1 4297 QDFFRBN $T=982700 578040 0 180 $X=970920 $Y=572620
X544 4284 4080 4273 2 1 4302 QDFFRBN $T=970920 598200 1 0 $X=970920 $Y=592780
X545 4297 4080 4273 2 1 4321 QDFFRBN $T=970920 598200 0 0 $X=970920 $Y=597820
X546 4299 585 4295 2 1 4353 QDFFRBN $T=971540 588120 1 0 $X=971540 $Y=582700
X547 4302 585 4295 2 1 4339 QDFFRBN $T=974020 588120 0 0 $X=974020 $Y=587740
X548 4283 585 619 2 1 622 QDFFRBN $T=977120 547800 1 0 $X=977120 $Y=542380
X549 4346 4080 4309 2 1 4317 QDFFRBN $T=990760 618360 1 180 $X=978980 $Y=617980
X550 4291 4080 4345 2 1 4366 QDFFRBN $T=980840 648600 0 0 $X=980840 $Y=648220
X551 4323 4080 4345 2 1 4328 QDFFRBN $T=981460 658680 1 0 $X=981460 $Y=653260
X552 4328 4080 4333 2 1 4360 QDFFRBN $T=981460 658680 0 0 $X=981460 $Y=658300
X553 4355 624 4333 2 1 4326 QDFFRBN $T=993240 678840 1 180 $X=981460 $Y=678460
X554 4331 4080 4313 2 1 4363 QDFFRBN $T=983320 638520 0 0 $X=983320 $Y=638140
X555 4339 585 4343 2 1 4372 QDFFRBN $T=986420 588120 0 0 $X=986420 $Y=587740
X556 4379 585 4330 2 1 4341 QDFFRBN $T=999440 557880 1 180 $X=987660 $Y=557500
X557 4354 4080 4313 2 1 4331 QDFFRBN $T=999440 638520 0 180 $X=987660 $Y=633100
X558 4384 585 4359 2 1 4348 QDFFRBN $T=1001300 547800 1 180 $X=989520 $Y=547420
X559 4348 585 4330 2 1 4379 QDFFRBN $T=989520 557880 1 0 $X=989520 $Y=552460
X560 4344 585 4343 2 1 4388 QDFFRBN $T=989520 578040 1 0 $X=989520 $Y=572620
X561 4353 585 4343 2 1 4380 QDFFRBN $T=989520 588120 1 0 $X=989520 $Y=582700
X562 4385 4080 4367 2 1 4357 QDFFRBN $T=1003780 628440 1 180 $X=992000 $Y=628060
X563 4363 4080 4345 2 1 4404 QDFFRBN $T=993860 648600 1 0 $X=993860 $Y=643180
X564 4366 4080 4333 2 1 4405 QDFFRBN $T=993860 648600 0 0 $X=993860 $Y=648220
X565 4360 4080 4333 2 1 4365 QDFFRBN $T=1006260 658680 1 180 $X=994480 $Y=658300
X566 4391 4080 4333 2 1 4362 QDFFRBN $T=1006260 668760 0 180 $X=994480 $Y=663340
X567 4368 624 4387 2 1 4396 QDFFRBN $T=994480 678840 1 0 $X=994480 $Y=673420
X568 4372 585 4343 2 1 4420 QDFFRBN $T=1001920 588120 1 0 $X=1001920 $Y=582700
X569 639 585 4359 2 1 4386 QDFFRBN $T=1014320 547800 1 180 $X=1002540 $Y=547420
X570 4388 585 4409 2 1 4389 QDFFRBN $T=1002540 567960 0 0 $X=1002540 $Y=567580
X571 4389 585 4343 2 1 4423 QDFFRBN $T=1002540 578040 1 0 $X=1002540 $Y=572620
X572 4390 624 4407 2 1 4416 QDFFRBN $T=1002540 699000 0 0 $X=1002540 $Y=698620
X573 4415 585 637 2 1 4384 QDFFRBN $T=1014940 557880 0 180 $X=1003160 $Y=552460
X574 4386 585 4409 2 1 4415 QDFFRBN $T=1003160 567960 1 0 $X=1003160 $Y=562540
X575 4426 4080 4367 2 1 4385 QDFFRBN $T=1015560 628440 1 180 $X=1003780 $Y=628060
X576 4401 624 641 2 1 643 QDFFRBN $T=1005640 719160 1 0 $X=1005640 $Y=713740
X577 4402 4080 4345 2 1 4426 QDFFRBN $T=1006260 638520 1 0 $X=1006260 $Y=633100
X578 642 624 4407 2 1 4390 QDFFRBN $T=1018040 709080 0 180 $X=1006260 $Y=703660
X579 4404 4080 4345 2 1 4432 QDFFRBN $T=1006880 648600 1 0 $X=1006880 $Y=643180
X580 4405 4080 4418 2 1 4419 QDFFRBN $T=1006880 648600 0 0 $X=1006880 $Y=648220
X581 4425 4080 4410 2 1 4403 QDFFRBN $T=1019280 608280 0 180 $X=1007500 $Y=602860
X582 4403 4080 4410 2 1 4408 QDFFRBN $T=1008740 608280 0 0 $X=1008740 $Y=607900
X583 4411 4080 4428 2 1 4441 QDFFRBN $T=1011220 598200 1 0 $X=1011220 $Y=592780
X584 4380 4080 4428 2 1 4444 QDFFRBN $T=1011840 588120 0 0 $X=1011840 $Y=587740
X585 4412 4080 4410 2 1 4440 QDFFRBN $T=1011840 618360 1 0 $X=1011840 $Y=612940
X586 4413 624 4387 2 1 4414 QDFFRBN $T=1012460 668760 0 0 $X=1012460 $Y=668380
X587 4414 624 4387 2 1 4443 QDFFRBN $T=1012460 678840 1 0 $X=1012460 $Y=673420
X588 4442 624 4387 2 1 4413 QDFFRBN $T=1024860 668760 0 180 $X=1013080 $Y=663340
X589 4419 4080 4418 2 1 4442 QDFFRBN $T=1014320 658680 1 0 $X=1014320 $Y=653260
X590 4420 585 4428 2 1 4411 QDFFRBN $T=1014940 588120 1 0 $X=1014940 $Y=582700
X591 4445 585 644 2 1 4417 QDFFRBN $T=1027340 547800 0 180 $X=1015560 $Y=542380
X592 4423 585 4428 2 1 4447 QDFFRBN $T=1015560 578040 1 0 $X=1015560 $Y=572620
X593 4421 585 4409 2 1 4448 QDFFRBN $T=1016180 547800 0 0 $X=1016180 $Y=547420
X594 4446 585 4409 2 1 4421 QDFFRBN $T=1027960 557880 1 180 $X=1016180 $Y=557500
X595 4447 585 4427 2 1 4422 QDFFRBN $T=1027960 567960 1 180 $X=1016180 $Y=567580
X596 4431 4080 4437 2 1 4402 QDFFRBN $T=1030440 628440 0 180 $X=1018660 $Y=623020
X597 4430 624 4406 2 1 4459 QDFFRBN $T=1018660 688920 0 0 $X=1018660 $Y=688540
X598 4456 4451 4438 2 1 4429 QDFFRBN $T=1031060 608280 0 180 $X=1019280 $Y=602860
X599 4461 624 641 2 1 4401 QDFFRBN $T=1031060 719160 0 180 $X=1019280 $Y=713740
X600 4458 4080 4418 2 1 4433 QDFFRBN $T=1032300 648600 1 180 $X=1020520 $Y=648220
X601 4434 624 4407 2 1 4435 QDFFRBN $T=1020520 699000 0 0 $X=1020520 $Y=698620
X602 4462 4451 4410 2 1 4439 QDFFRBN $T=1034780 608280 1 180 $X=1023000 $Y=607900
X603 4440 4451 4410 2 1 4436 QDFFRBN $T=1035400 618360 0 180 $X=1023620 $Y=612940
X604 4441 585 4438 2 1 4465 QDFFRBN $T=1024240 598200 1 0 $X=1024240 $Y=592780
X605 4444 585 4438 2 1 4470 QDFFRBN $T=1024860 588120 0 0 $X=1024860 $Y=587740
X606 4422 585 4427 2 1 4446 QDFFRBN $T=1025480 567960 1 0 $X=1025480 $Y=562540
X607 4443 624 4449 2 1 4477 QDFFRBN $T=1026720 668760 0 0 $X=1026720 $Y=668380
X608 4477 624 4449 2 1 4450 QDFFRBN $T=1039740 678840 0 180 $X=1027960 $Y=673420
X609 4448 585 4409 2 1 4453 QDFFRBN $T=1040360 547800 1 180 $X=1028580 $Y=547420
X610 4479 585 4409 2 1 4454 QDFFRBN $T=1040360 557880 1 180 $X=1028580 $Y=557500
X611 4453 585 4427 2 1 4485 QDFFRBN $T=1029200 567960 0 0 $X=1029200 $Y=567580
X612 4450 624 4449 2 1 4482 QDFFRBN $T=1029200 678840 0 0 $X=1029200 $Y=678460
X613 4429 4451 4438 2 1 4425 QDFFRBN $T=1042840 608280 0 180 $X=1031060 $Y=602860
X614 4459 624 4452 2 1 4497 QDFFRBN $T=1031060 688920 0 0 $X=1031060 $Y=688540
X615 649 624 641 2 1 4461 QDFFRBN $T=1045320 719160 0 180 $X=1033540 $Y=713740
X616 4463 624 4452 2 1 4488 QDFFRBN $T=1034160 709080 1 0 $X=1034160 $Y=703660
X617 4464 4451 4474 2 1 4457 QDFFRBN $T=1046560 638520 1 180 $X=1034780 $Y=638140
X618 4467 624 4452 2 1 4463 QDFFRBN $T=1046560 699000 1 180 $X=1034780 $Y=698620
X619 4488 624 4475 2 1 645 QDFFRBN $T=1046560 709080 1 180 $X=1034780 $Y=708700
X620 4493 624 4452 2 1 4467 QDFFRBN $T=1047180 699000 0 180 $X=1035400 $Y=693580
X621 4494 4451 4449 2 1 4468 QDFFRBN $T=1047800 668760 0 180 $X=1036020 $Y=663340
X622 4469 624 4487 2 1 4493 QDFFRBN $T=1036020 688920 1 0 $X=1036020 $Y=683500
X623 4499 4451 4438 2 1 4456 QDFFRBN $T=1048420 608280 1 180 $X=1036640 $Y=607900
X624 4495 4451 4437 2 1 4471 QDFFRBN $T=1048420 628440 0 180 $X=1036640 $Y=623020
X625 4465 650 4438 2 1 4472 QDFFRBN $T=1049040 588120 1 180 $X=1037260 $Y=587740
X626 4470 585 4490 2 1 4505 QDFFRBN $T=1037260 598200 1 0 $X=1037260 $Y=592780
X627 4472 585 4490 2 1 4498 QDFFRBN $T=1037880 588120 1 0 $X=1037880 $Y=582700
X628 4476 4451 4490 2 1 4499 QDFFRBN $T=1037880 618360 1 0 $X=1037880 $Y=612940
X629 4481 650 4484 2 1 4479 QDFFRBN $T=1051520 567960 0 180 $X=1039740 $Y=562540
X630 4468 4451 4449 2 1 4507 QDFFRBN $T=1040360 668760 0 0 $X=1040360 $Y=668380
X631 4482 624 4487 2 1 4469 QDFFRBN $T=1041600 678840 0 0 $X=1041600 $Y=678460
X632 4513 650 4484 2 1 4481 QDFFRBN $T=1054000 557880 1 180 $X=1042220 $Y=557500
X633 4485 585 4484 2 1 4489 QDFFRBN $T=1042220 567960 0 0 $X=1042220 $Y=567580
X634 4497 624 4487 2 1 4516 QDFFRBN $T=1046560 688920 0 0 $X=1046560 $Y=688540
X635 4498 650 4510 2 1 4506 QDFFRBN $T=1048420 578040 0 0 $X=1048420 $Y=577660
X636 4518 4451 4490 2 1 4476 QDFFRBN $T=1060820 608280 1 180 $X=1049040 $Y=607900
X637 4500 4451 4508 2 1 4520 QDFFRBN $T=1049040 648600 1 0 $X=1049040 $Y=643180
X638 4519 624 4475 2 1 4397 QDFFRBN $T=1060820 719160 0 180 $X=1049040 $Y=713740
X639 4505 650 4510 2 1 4525 QDFFRBN $T=1049660 598200 1 0 $X=1049660 $Y=592780
X640 4528 4451 4508 2 1 4496 QDFFRBN $T=1061440 638520 1 180 $X=1049660 $Y=638140
X641 4504 4451 4478 2 1 4500 QDFFRBN $T=1061440 658680 0 180 $X=1049660 $Y=653260
X642 4506 650 4490 2 1 4548 QDFFRBN $T=1050280 588120 0 0 $X=1050280 $Y=587740
X643 4522 4451 4510 2 1 4502 QDFFRBN $T=1062060 598200 1 180 $X=1050280 $Y=597820
X644 4502 4451 4510 2 1 4518 QDFFRBN $T=1050280 608280 1 0 $X=1050280 $Y=602860
X645 4533 4451 4478 2 1 4504 QDFFRBN $T=1062060 658680 1 180 $X=1050280 $Y=658300
X646 4507 4451 4449 2 1 4531 QDFFRBN $T=1050280 668760 1 0 $X=1050280 $Y=663340
X647 652 650 4523 2 1 4511 QDFFRBN $T=1052760 547800 1 0 $X=1052760 $Y=542380
X648 4511 650 4523 2 1 4544 QDFFRBN $T=1053380 547800 0 0 $X=1053380 $Y=547420
X649 4531 4451 4514 2 1 4512 QDFFRBN $T=1065780 668760 1 180 $X=1054000 $Y=668380
X650 4489 650 4484 2 1 4542 QDFFRBN $T=1055240 557880 1 0 $X=1055240 $Y=552460
X651 4512 624 4487 2 1 4547 QDFFRBN $T=1055240 678840 0 0 $X=1055240 $Y=678460
X652 4543 650 4484 2 1 4513 QDFFRBN $T=1067640 557880 1 180 $X=1055860 $Y=557500
X653 4538 624 4475 2 1 654 QDFFRBN $T=1068880 709080 1 180 $X=1057100 $Y=708700
X654 4515 4451 4508 2 1 4555 QDFFRBN $T=1057720 638520 1 0 $X=1057720 $Y=633100
X655 4525 650 4532 2 1 4546 QDFFRBN $T=1061440 588120 1 0 $X=1061440 $Y=582700
X656 4548 650 4510 2 1 4522 QDFFRBN $T=1073840 598200 0 180 $X=1062060 $Y=592780
X657 4553 4451 4534 2 1 4526 QDFFRBN $T=1073840 608280 1 180 $X=1062060 $Y=607900
X658 4549 624 4475 2 1 4527 QDFFRBN $T=1073840 709080 0 180 $X=1062060 $Y=703660
X659 4527 624 653 2 1 4519 QDFFRBN $T=1062060 719160 1 0 $X=1062060 $Y=713740
X660 4530 4451 4534 2 1 4554 QDFFRBN $T=1063300 628440 1 0 $X=1063300 $Y=623020
X661 4552 4451 4536 2 1 4528 QDFFRBN $T=1075080 638520 1 180 $X=1063300 $Y=638140
X662 4529 4451 4541 2 1 4552 QDFFRBN $T=1063300 648600 1 0 $X=1063300 $Y=643180
X663 4561 4451 4541 2 1 4535 QDFFRBN $T=1076940 658680 0 180 $X=1065160 $Y=653260
X664 4535 4451 4541 2 1 4533 QDFFRBN $T=1076940 658680 1 180 $X=1065160 $Y=658300
X665 4540 624 4514 2 1 4567 QDFFRBN $T=1067640 678840 1 0 $X=1067640 $Y=673420
X666 4544 650 4523 2 1 4545 QDFFRBN $T=1068260 547800 0 0 $X=1068260 $Y=547420
X667 4542 650 4523 2 1 4572 QDFFRBN $T=1068260 557880 0 0 $X=1068260 $Y=557500
X668 4545 650 656 2 1 657 QDFFRBN $T=1069500 547800 1 0 $X=1069500 $Y=542380
X669 4554 4451 4534 2 1 4565 QDFFRBN $T=1073840 628440 0 0 $X=1073840 $Y=628060
X670 4573 4451 4551 2 1 4553 QDFFRBN $T=1086240 608280 1 180 $X=1074460 $Y=607900
X671 4574 624 4514 2 1 4540 QDFFRBN $T=1086240 678840 1 180 $X=1074460 $Y=678460
X672 4557 624 4566 2 1 4574 QDFFRBN $T=1074460 688920 1 0 $X=1074460 $Y=683500
X673 4577 624 4566 2 1 4556 QDFFRBN $T=1086240 699000 0 180 $X=1074460 $Y=693580
X674 4556 624 4566 2 1 4557 QDFFRBN $T=1086240 699000 1 180 $X=1074460 $Y=698620
X675 4563 650 4569 2 1 4564 QDFFRBN $T=1075080 578040 1 0 $X=1075080 $Y=572620
X676 4559 4451 4551 2 1 4573 QDFFRBN $T=1075080 608280 1 0 $X=1075080 $Y=602860
X677 4582 650 4569 2 1 4543 QDFFRBN $T=1087480 567960 1 180 $X=1075700 $Y=567580
X678 4564 650 4568 2 1 4588 QDFFRBN $T=1075700 578040 0 0 $X=1075700 $Y=577660
X679 4565 4451 4536 2 1 4589 QDFFRBN $T=1075700 638520 1 0 $X=1075700 $Y=633100
X680 4555 4451 4536 2 1 4592 QDFFRBN $T=1076320 638520 0 0 $X=1076320 $Y=638140
X681 4583 4451 4536 2 1 4529 QDFFRBN $T=1088100 648600 0 180 $X=1076320 $Y=643180
X682 4595 650 656 2 1 4571 QDFFRBN $T=1093680 547800 1 180 $X=1081900 $Y=547420
X683 4572 650 4569 2 1 4596 QDFFRBN $T=1081900 557880 0 0 $X=1081900 $Y=557500
X684 4571 650 658 2 1 659 QDFFRBN $T=1082520 547800 1 0 $X=1082520 $Y=542380
X685 4608 4451 4551 2 1 4576 QDFFRBN $T=1098640 618360 0 180 $X=1086860 $Y=612940
X686 4602 4451 4591 2 1 4579 QDFFRBN $T=1099260 608280 1 180 $X=1087480 $Y=607900
X687 4576 4451 4591 2 1 4606 QDFFRBN $T=1087480 618360 0 0 $X=1087480 $Y=617980
X688 4580 4451 4597 2 1 4560 QDFFRBN $T=1088100 598200 1 0 $X=1088100 $Y=592780
X689 4581 624 4566 2 1 4577 QDFFRBN $T=1099880 699000 0 180 $X=1088100 $Y=693580
X690 4588 650 4568 2 1 4605 QDFFRBN $T=1089340 578040 0 0 $X=1089340 $Y=577660
X691 4605 650 4568 2 1 4585 QDFFRBN $T=1101120 588120 0 180 $X=1089340 $Y=582700
X692 4585 650 4568 2 1 4580 QDFFRBN $T=1101120 588120 1 180 $X=1089340 $Y=587740
X693 4589 4451 4600 2 1 4593 QDFFRBN $T=1089340 638520 1 0 $X=1089340 $Y=633100
X694 4587 4451 4594 2 1 4612 QDFFRBN $T=1089340 658680 1 0 $X=1089340 $Y=653260
X695 4610 624 4562 2 1 4586 QDFFRBN $T=1101120 668760 1 180 $X=1089340 $Y=668380
X696 4592 4451 4600 2 1 4587 QDFFRBN $T=1089960 638520 0 0 $X=1089960 $Y=638140
X697 4593 4451 4600 2 1 4621 QDFFRBN $T=1091200 628440 0 0 $X=1091200 $Y=628060
X698 4596 650 4601 2 1 4614 QDFFRBN $T=1094920 557880 0 0 $X=1094920 $Y=557500
X699 661 650 658 2 1 4595 QDFFRBN $T=1107320 547800 1 180 $X=1095540 $Y=547420
X700 4579 4451 4597 2 1 4617 QDFFRBN $T=1095540 608280 1 0 $X=1095540 $Y=602860
X701 660 650 658 2 1 4619 QDFFRBN $T=1096160 547800 1 0 $X=1096160 $Y=542380
X702 4616 650 4604 2 1 4582 QDFFRBN $T=1107940 567960 1 180 $X=1096160 $Y=567580
X703 4598 650 4601 2 1 4616 QDFFRBN $T=1096160 578040 1 0 $X=1096160 $Y=572620
X704 4617 650 4597 2 1 4599 QDFFRBN $T=1108560 598200 1 180 $X=1096780 $Y=597820
X705 4625 4451 4591 2 1 4608 QDFFRBN $T=1112280 608280 1 180 $X=1100500 $Y=607900
X706 4606 4451 4591 2 1 4602 QDFFRBN $T=1112280 618360 1 180 $X=1100500 $Y=617980
X707 4599 650 4613 2 1 4623 QDFFRBN $T=1101120 598200 1 0 $X=1101120 $Y=592780
X708 4624 4451 4562 2 1 4610 QDFFRBN $T=1114140 668760 1 180 $X=1102360 $Y=668380
X709 4611 624 4562 2 1 4624 QDFFRBN $T=1102980 668760 1 0 $X=1102980 $Y=663340
X710 4628 4451 4594 2 1 4590 QDFFRBN $T=1116000 648600 1 180 $X=1104220 $Y=648220
X711 4614 650 4601 2 1 4622 QDFFRBN $T=1105460 567960 1 0 $X=1105460 $Y=562540
X712 4615 4451 4600 2 1 4628 QDFFRBN $T=1105460 638520 0 0 $X=1105460 $Y=638140
X713 4619 650 658 2 1 4634 QDFFRBN $T=1108560 547800 0 0 $X=1108560 $Y=547420
X714 4621 4451 4618 2 1 4629 QDFFRBN $T=1109180 628440 0 0 $X=1109180 $Y=628060
X715 4622 650 4604 2 1 4630 QDFFRBN $T=1109800 567960 0 0 $X=1109800 $Y=567580
X716 4631 650 4601 2 1 4598 QDFFRBN $T=1121580 578040 0 180 $X=1109800 $Y=572620
X717 4629 4451 4618 2 1 4615 QDFFRBN $T=1121580 638520 0 180 $X=1109800 $Y=633100
X718 4630 650 4604 2 1 4620 QDFFRBN $T=1122200 578040 1 180 $X=1110420 $Y=577660
X719 4623 650 4613 2 1 4631 QDFFRBN $T=1110420 588120 1 0 $X=1110420 $Y=582700
X720 4620 650 4613 2 1 4633 QDFFRBN $T=1113520 588120 0 0 $X=1113520 $Y=587740
X721 4632 4451 4618 2 1 4625 QDFFRBN $T=1125300 608280 1 180 $X=1113520 $Y=607900
X722 4633 4451 4613 2 1 4627 QDFFRBN $T=1125920 598200 0 180 $X=1114140 $Y=592780
X723 4627 4451 4618 2 1 4632 QDFFRBN $T=1114140 608280 1 0 $X=1114140 $Y=602860
X724 4634 650 663 2 1 662 QDFFRBN $T=1127780 547800 0 180 $X=1116000 $Y=542380
X725 683 2 704 1 INV1S $T=264740 608280 1 0 $X=264740 $Y=602860
X726 692 2 718 1 INV1S $T=265360 578040 1 0 $X=265360 $Y=572620
X727 713 2 725 1 INV1S $T=269700 618360 1 0 $X=269700 $Y=612940
X728 718 2 701 1 INV1S $T=272180 567960 0 0 $X=272180 $Y=567580
X729 705 2 735 1 INV1S $T=276520 588120 0 0 $X=276520 $Y=587740
X730 727 2 753 1 INV1S $T=283340 628440 0 180 $X=282100 $Y=623020
X731 684 2 760 1 INV1S $T=285820 608280 1 0 $X=285820 $Y=602860
X732 702 2 755 1 INV1S $T=288300 628440 1 180 $X=287060 $Y=628060
X733 769 2 757 1 INV1S $T=288920 567960 1 180 $X=287680 $Y=567580
X734 782 2 785 1 INV1S $T=288920 588120 0 0 $X=288920 $Y=587740
X735 789 2 780 1 INV1S $T=291400 668760 1 180 $X=290160 $Y=668380
X736 839 2 810 1 INV1S $T=295120 699000 0 180 $X=293880 $Y=693580
X737 813 2 824 1 INV1S $T=295120 608280 0 0 $X=295120 $Y=607900
X738 823 2 818 1 INV1S $T=296360 658680 0 180 $X=295120 $Y=653260
X739 772 2 826 1 INV1S $T=295740 598200 1 0 $X=295740 $Y=592780
X740 830 2 836 1 INV1S $T=296980 598200 1 0 $X=296980 $Y=592780
X741 827 2 825 1 INV1S $T=298840 648600 1 180 $X=297600 $Y=648220
X742 856 2 849 1 INV1S $T=302560 648600 0 180 $X=301320 $Y=643180
X743 840 2 860 1 INV1S $T=301940 598200 0 0 $X=301940 $Y=597820
X744 844 2 863 1 INV1S $T=303180 658680 1 0 $X=303180 $Y=653260
X745 847 2 873 1 INV1S $T=304420 598200 1 0 $X=304420 $Y=592780
X746 891 2 870 1 INV1S $T=306900 638520 0 180 $X=305660 $Y=633100
X747 787 2 890 1 INV1S $T=307520 618360 1 0 $X=307520 $Y=612940
X748 892 2 881 1 INV1S $T=308760 678840 0 180 $X=307520 $Y=673420
X749 16 2 898 1 INV1S $T=308760 547800 1 0 $X=308760 $Y=542380
X750 872 2 879 1 INV1S $T=310000 648600 0 180 $X=308760 $Y=643180
X751 875 2 883 1 INV1S $T=310620 658680 0 180 $X=309380 $Y=653260
X752 852 2 887 1 INV1S $T=310620 658680 1 180 $X=309380 $Y=658300
X753 799 2 929 1 INV1S $T=316820 628440 1 180 $X=315580 $Y=628060
X754 934 2 920 1 INV1S $T=316820 638520 0 180 $X=315580 $Y=633100
X755 876 2 911 1 INV1S $T=317440 658680 1 180 $X=316200 $Y=658300
X756 900 2 951 1 INV1S $T=316820 557880 1 0 $X=316820 $Y=552460
X757 950 2 869 1 INV1S $T=318680 648600 1 180 $X=317440 $Y=648220
X758 945 2 921 1 INV1S $T=319300 658680 1 180 $X=318060 $Y=658300
X759 21 2 956 1 INV1S $T=319300 547800 0 0 $X=319300 $Y=547420
X760 894 2 930 1 INV1S $T=321160 608280 1 180 $X=319920 $Y=607900
X761 962 2 937 1 INV1S $T=321160 668760 1 180 $X=319920 $Y=668380
X762 22 2 965 1 INV1S $T=320540 547800 0 0 $X=320540 $Y=547420
X763 964 2 972 1 INV1S $T=324260 688920 0 180 $X=323020 $Y=683500
X764 996 2 992 1 INV1S $T=329220 608280 0 180 $X=327980 $Y=602860
X765 923 2 1026 1 INV1S $T=329840 557880 1 0 $X=329840 $Y=552460
X766 927 2 1002 1 INV1S $T=329840 638520 1 0 $X=329840 $Y=633100
X767 960 2 988 1 INV1S $T=330460 588120 0 0 $X=330460 $Y=587740
X768 966 2 991 1 INV1S $T=331080 588120 1 0 $X=331080 $Y=582700
X769 31 2 1048 1 INV1S $T=335420 547800 1 0 $X=335420 $Y=542380
X770 1037 2 1046 1 INV1S $T=337280 648600 1 180 $X=336040 $Y=648220
X771 963 2 1025 1 INV1S $T=337280 668760 0 180 $X=336040 $Y=663340
X772 1058 2 1012 1 INV1S $T=338520 678840 0 180 $X=337280 $Y=673420
X773 1042 2 1013 1 INV1S $T=337900 598200 0 0 $X=337900 $Y=597820
X774 40 2 1063 1 INV1S $T=339140 547800 1 0 $X=339140 $Y=542380
X775 1067 2 1076 1 INV1S $T=340380 688920 1 0 $X=340380 $Y=683500
X776 1065 2 1047 1 INV1S $T=341620 658680 1 0 $X=341620 $Y=653260
X777 1045 2 1077 1 INV1S $T=342240 628440 0 0 $X=342240 $Y=628060
X778 42 2 1087 1 INV1S $T=342240 719160 1 0 $X=342240 $Y=713740
X779 1082 2 1057 1 INV1S $T=344720 598200 1 180 $X=343480 $Y=597820
X780 1066 2 1022 1 INV1S $T=345340 658680 0 0 $X=345340 $Y=658300
X781 946 2 1106 1 INV1S $T=347200 618360 0 0 $X=347200 $Y=617980
X782 1116 2 1020 1 INV1S $T=348440 638520 0 180 $X=347200 $Y=633100
X783 1117 2 1101 1 INV1S $T=349060 608280 0 180 $X=347820 $Y=602860
X784 1111 2 1094 1 INV1S $T=349060 608280 1 180 $X=347820 $Y=607900
X785 1098 2 1055 1 INV1S $T=349060 668760 1 180 $X=347820 $Y=668380
X786 1079 2 1112 1 INV1S $T=347820 709080 0 0 $X=347820 $Y=708700
X787 50 2 1061 1 INV1S $T=350920 658680 0 180 $X=349680 $Y=653260
X788 954 2 1119 1 INV1S $T=350920 567960 0 0 $X=350920 $Y=567580
X789 1160 2 1124 1 INV1S $T=353400 648600 1 180 $X=352160 $Y=648220
X790 1139 2 1136 1 INV1S $T=354020 628440 0 180 $X=352780 $Y=623020
X791 1133 2 1143 1 INV1S $T=355880 578040 1 180 $X=354640 $Y=577660
X792 1125 2 1166 1 INV1S $T=357740 578040 0 0 $X=357740 $Y=577660
X793 1156 2 1162 1 INV1S $T=360220 567960 0 180 $X=358980 $Y=562540
X794 1176 2 1163 1 INV1S $T=360220 608280 0 180 $X=358980 $Y=602860
X795 1097 2 1175 1 INV1S $T=359600 618360 1 0 $X=359600 $Y=612940
X796 1065 2 1185 1 INV1S $T=360220 638520 1 0 $X=360220 $Y=633100
X797 1155 2 1179 1 INV1S $T=360220 648600 1 0 $X=360220 $Y=643180
X798 1211 2 868 1 INV1S $T=362080 648600 1 180 $X=360840 $Y=648220
X799 1085 2 1194 1 INV1S $T=362080 567960 0 0 $X=362080 $Y=567580
X800 1044 2 1210 1 INV1S $T=362700 557880 0 0 $X=362700 $Y=557500
X801 1158 2 1184 1 INV1S $T=364560 578040 1 180 $X=363320 $Y=577660
X802 1172 2 1208 1 INV1S $T=364560 567960 1 0 $X=364560 $Y=562540
X803 1126 2 1226 1 INV1S $T=366420 557880 0 0 $X=366420 $Y=557500
X804 1219 2 1224 1 INV1S $T=366420 588120 0 0 $X=366420 $Y=587740
X805 1227 2 1200 1 INV1S $T=368280 618360 0 180 $X=367040 $Y=612940
X806 1211 2 950 1 INV1S $T=367040 648600 0 0 $X=367040 $Y=648220
X807 1217 2 1157 1 INV1S $T=367660 719160 1 0 $X=367660 $Y=713740
X808 1167 2 1229 1 INV1S $T=368280 557880 1 0 $X=368280 $Y=552460
X809 1215 2 1231 1 INV1S $T=368280 618360 1 0 $X=368280 $Y=612940
X810 1144 2 1222 1 INV1S $T=368280 699000 1 0 $X=368280 $Y=693580
X811 1220 2 1256 1 INV1S $T=370760 557880 1 0 $X=370760 $Y=552460
X812 1247 2 1180 1 INV1S $T=370760 618360 0 0 $X=370760 $Y=617980
X813 1181 2 1242 1 INV1S $T=372620 699000 0 180 $X=371380 $Y=693580
X814 1132 2 1245 1 INV1S $T=373860 557880 1 180 $X=372620 $Y=557500
X815 1259 2 1243 1 INV1S $T=373860 608280 0 180 $X=372620 $Y=602860
X816 1264 2 1258 1 INV1S $T=373860 638520 0 180 $X=372620 $Y=633100
X817 1263 2 1233 1 INV1S $T=374480 588120 1 180 $X=373240 $Y=587740
X818 1141 2 1260 1 INV1S $T=373860 688920 0 0 $X=373860 $Y=688540
X819 60 2 1277 1 INV1S $T=375100 719160 1 0 $X=375100 $Y=713740
X820 1280 2 1255 1 INV1S $T=376960 618360 0 180 $X=375720 $Y=612940
X821 1145 2 1273 1 INV1S $T=377580 547800 0 0 $X=377580 $Y=547420
X822 1300 2 1296 1 INV1S $T=380060 648600 0 0 $X=380060 $Y=648220
X823 1309 2 1298 1 INV1S $T=381920 628440 0 180 $X=380680 $Y=623020
X824 1319 2 1352 1 INV1S $T=386260 547800 0 0 $X=386260 $Y=547420
X825 1336 2 1345 1 INV1S $T=387500 547800 1 0 $X=387500 $Y=542380
X826 1223 2 1228 1 INV1S $T=390600 638520 0 0 $X=390600 $Y=638140
X827 1339 2 1201 1 INV1S $T=391220 628440 1 0 $X=391220 $Y=623020
X828 74 2 1083 1 INV1S $T=393700 688920 0 180 $X=392460 $Y=683500
X829 1371 2 1365 1 INV1S $T=394320 618360 1 180 $X=393080 $Y=617980
X830 1381 2 1291 1 INV1S $T=396180 658680 0 180 $X=394940 $Y=653260
X831 74 2 985 1 INV1S $T=396800 567960 1 180 $X=395560 $Y=567580
X832 1391 2 1267 1 INV1S $T=398040 648600 1 180 $X=396800 $Y=648220
X833 1381 2 1391 1 INV1S $T=396800 658680 1 0 $X=396800 $Y=653260
X834 1355 2 1375 1 INV1S $T=398660 598200 0 180 $X=397420 $Y=592780
X835 1387 2 1386 1 INV1S $T=399280 709080 0 180 $X=398040 $Y=703660
X836 1406 2 1408 1 INV1S $T=399900 618360 0 0 $X=399900 $Y=617980
X837 1394 2 77 1 INV1S $T=401140 719160 0 180 $X=399900 $Y=713740
X838 78 2 1393 1 INV1S $T=402380 699000 1 180 $X=401140 $Y=698620
X839 1369 2 1421 1 INV1S $T=402380 658680 1 0 $X=402380 $Y=653260
X840 1400 2 1406 1 INV1S $T=403000 618360 1 0 $X=403000 $Y=612940
X841 74 2 1415 1 INV1S $T=404240 578040 0 0 $X=404240 $Y=577660
X842 1383 2 1431 1 INV1S $T=405480 567960 1 0 $X=405480 $Y=562540
X843 1436 2 1417 1 INV1S $T=406720 648600 1 0 $X=406720 $Y=643180
X844 87 2 1414 1 INV1S $T=409200 547800 0 180 $X=407960 $Y=542380
X845 1465 2 1430 1 INV1S $T=409200 688920 0 180 $X=407960 $Y=683500
X846 1425 2 1458 1 INV1S $T=410440 578040 0 0 $X=410440 $Y=577660
X847 1455 2 1396 1 INV1S $T=411680 588120 0 180 $X=410440 $Y=582700
X848 1471 2 1381 1 INV1S $T=412300 648600 1 180 $X=411060 $Y=648220
X849 1461 2 1459 1 INV1S $T=413540 618360 0 180 $X=412300 $Y=612940
X850 1460 2 1477 1 INV1S $T=413540 598200 0 0 $X=413540 $Y=597820
X851 96 2 1446 1 INV1S $T=415400 547800 0 180 $X=414160 $Y=542380
X852 1468 2 92 1 INV1S $T=416020 719160 0 180 $X=414780 $Y=713740
X853 1457 2 1495 1 INV1S $T=416020 567960 1 0 $X=416020 $Y=562540
X854 1484 2 1447 1 INV1S $T=417260 638520 0 180 $X=416020 $Y=633100
X855 1491 2 1490 1 INV1S $T=417260 588120 1 0 $X=417260 $Y=582700
X856 1211 2 1497 1 INV1S $T=417260 648600 1 0 $X=417260 $Y=643180
X857 1466 2 1496 1 INV1S $T=420360 608280 0 180 $X=419120 $Y=602860
X858 1467 2 1505 1 INV1S $T=419740 678840 1 0 $X=419740 $Y=673420
X859 1508 2 1515 1 INV1S $T=420980 598200 1 0 $X=420980 $Y=592780
X860 1504 2 1527 1 INV1S $T=424080 648600 0 0 $X=424080 $Y=648220
X861 1529 2 1511 1 INV1S $T=425320 578040 0 0 $X=425320 $Y=577660
X862 1315 2 1499 1 INV1S $T=425940 638520 1 0 $X=425940 $Y=633100
X863 1539 2 1500 1 INV1S $T=427180 688920 1 180 $X=425940 $Y=688540
X864 1462 2 1520 1 INV1S $T=426560 578040 0 0 $X=426560 $Y=577660
X865 1533 2 1517 1 INV1S $T=428420 547800 0 180 $X=427180 $Y=542380
X866 1541 2 1530 1 INV1S $T=428420 638520 0 180 $X=427180 $Y=633100
X867 1211 2 1542 1 INV1S $T=427180 648600 1 0 $X=427180 $Y=643180
X868 1547 2 1552 1 INV1S $T=429660 688920 1 0 $X=429660 $Y=683500
X869 1521 2 1563 1 INV1S $T=431520 608280 1 0 $X=431520 $Y=602860
X870 1548 2 1560 1 INV1S $T=431520 618360 1 0 $X=431520 $Y=612940
X871 1575 2 1553 1 INV1S $T=434620 567960 1 180 $X=433380 $Y=567580
X872 1571 2 1582 1 INV1S $T=434620 608280 0 0 $X=434620 $Y=607900
X873 1557 2 1580 1 INV1S $T=435240 699000 1 0 $X=435240 $Y=693580
X874 1586 2 1576 1 INV1S $T=437720 567960 0 180 $X=436480 $Y=562540
X875 1433 2 1587 1 INV1S $T=436480 638520 0 0 $X=436480 $Y=638140
X876 1574 2 1564 1 INV1S $T=437100 618360 1 0 $X=437100 $Y=612940
X877 1589 2 1559 1 INV1S $T=438340 688920 0 180 $X=437100 $Y=683500
X878 1598 2 1584 1 INV1S $T=440820 709080 0 180 $X=439580 $Y=703660
X879 1599 2 1593 1 INV1S $T=441440 668760 1 180 $X=440200 $Y=668380
X880 1554 2 1603 1 INV1S $T=440820 578040 1 0 $X=440820 $Y=572620
X881 1579 2 1615 1 INV1S $T=441440 618360 0 0 $X=441440 $Y=617980
X882 1592 2 1618 1 INV1S $T=442680 567960 0 0 $X=442680 $Y=567580
X883 1526 2 1622 1 INV1S $T=442680 618360 0 0 $X=442680 $Y=617980
X884 1600 2 1640 1 INV1S $T=447020 618360 0 0 $X=447020 $Y=617980
X885 1627 2 1648 1 INV1S $T=449500 628440 0 0 $X=449500 $Y=628060
X886 1651 2 1646 1 INV1S $T=450740 699000 0 180 $X=449500 $Y=693580
X887 1606 2 1638 1 INV1S $T=450120 578040 1 0 $X=450120 $Y=572620
X888 1394 2 125 1 INV1S $T=450740 709080 0 0 $X=450740 $Y=708700
X889 1597 2 1661 1 INV1S $T=451980 567960 1 0 $X=451980 $Y=562540
X890 1608 2 1631 1 INV1S $T=453220 638520 1 180 $X=451980 $Y=638140
X891 1649 2 1658 1 INV1S $T=453220 699000 0 180 $X=451980 $Y=693580
X892 1642 2 1662 1 INV1S $T=452600 638520 1 0 $X=452600 $Y=633100
X893 1664 2 1666 1 INV1S $T=453840 709080 1 0 $X=453840 $Y=703660
X894 1671 2 1647 1 INV1S $T=455700 688920 1 180 $X=454460 $Y=688540
X895 1689 2 1688 1 INV1S $T=458800 578040 1 0 $X=458800 $Y=572620
X896 1693 2 1660 1 INV1S $T=460660 547800 0 0 $X=460660 $Y=547420
X897 1678 2 1703 1 INV1S $T=460660 709080 0 0 $X=460660 $Y=708700
X898 74 2 1699 1 INV1S $T=462520 638520 0 0 $X=462520 $Y=638140
X899 1675 2 1704 1 INV1S $T=463760 699000 0 0 $X=463760 $Y=698620
X900 1686 2 1717 1 INV1S $T=465620 547800 0 0 $X=465620 $Y=547420
X901 141 2 1728 1 INV1S $T=466240 719160 1 0 $X=466240 $Y=713740
X902 1749 2 1751 1 INV1S $T=469960 618360 1 0 $X=469960 $Y=612940
X903 1738 2 1759 1 INV1S $T=470580 567960 1 0 $X=470580 $Y=562540
X904 1719 2 1747 1 INV1S $T=470580 709080 0 0 $X=470580 $Y=708700
X905 1665 2 1770 1 INV1S $T=472440 648600 1 0 $X=472440 $Y=643180
X906 1713 2 1765 1 INV1S $T=474300 578040 0 180 $X=473060 $Y=572620
X907 1776 2 1758 1 INV1S $T=475540 618360 1 180 $X=474300 $Y=617980
X908 1772 2 1780 1 INV1S $T=474920 567960 1 0 $X=474920 $Y=562540
X909 1773 2 1799 1 INV1S $T=475540 578040 1 0 $X=475540 $Y=572620
X910 1774 2 1784 1 INV1S $T=475540 598200 1 0 $X=475540 $Y=592780
X911 1752 2 1787 1 INV1S $T=475540 648600 1 0 $X=475540 $Y=643180
X912 1741 2 1788 1 INV1S $T=475540 658680 1 0 $X=475540 $Y=653260
X913 1745 2 154 1 INV1S $T=476160 668760 0 0 $X=476160 $Y=668380
X914 1742 2 1778 1 INV1S $T=476160 688920 1 0 $X=476160 $Y=683500
X915 1781 2 1790 1 INV1S $T=476780 608280 1 0 $X=476780 $Y=602860
X916 1746 2 1783 1 INV1S $T=477400 567960 0 0 $X=477400 $Y=567580
X917 1777 2 1812 1 INV1S $T=477400 588120 1 0 $X=477400 $Y=582700
X918 1743 2 1793 1 INV1S $T=477400 598200 1 0 $X=477400 $Y=592780
X919 1736 2 1782 1 INV1S $T=478640 608280 1 180 $X=477400 $Y=607900
X920 1748 2 1829 1 INV1S $T=481740 578040 0 0 $X=481740 $Y=577660
X921 1750 2 155 1 INV1S $T=481740 678840 1 0 $X=481740 $Y=673420
X922 1779 2 156 1 INV1S $T=482360 699000 0 0 $X=482360 $Y=698620
X923 1828 2 157 1 INV1S $T=483600 709080 0 0 $X=483600 $Y=708700
X924 1731 2 1840 1 INV1S $T=486080 557880 1 0 $X=486080 $Y=552460
X925 1824 2 162 1 INV1S $T=488560 638520 0 0 $X=488560 $Y=638140
X926 1825 2 1856 1 INV1S $T=488560 668760 1 0 $X=488560 $Y=663340
X927 1836 2 1864 1 INV1S $T=490420 608280 0 0 $X=490420 $Y=607900
X928 1859 2 159 1 INV1S $T=491040 688920 0 0 $X=491040 $Y=688540
X929 1870 2 1877 1 INV1S $T=493520 567960 0 0 $X=493520 $Y=567580
X930 1874 2 1843 1 INV1S $T=493520 628440 0 0 $X=493520 $Y=628060
X931 1873 2 1868 1 INV1S $T=494140 618360 0 0 $X=494140 $Y=617980
X932 1855 2 1879 1 INV1S $T=494140 658680 0 0 $X=494140 $Y=658300
X933 1882 2 1860 1 INV1S $T=494760 608280 0 0 $X=494760 $Y=607900
X934 1884 2 1823 1 INV1S $T=496620 557880 0 180 $X=495380 $Y=552460
X935 1887 2 1853 1 INV1S $T=496000 588120 1 0 $X=496000 $Y=582700
X936 1869 2 1889 1 INV1S $T=496000 678840 0 0 $X=496000 $Y=678460
X937 1892 2 1835 1 INV1S $T=499720 557880 1 180 $X=498480 $Y=557500
X938 1900 2 1875 1 INV1S $T=499100 578040 0 0 $X=499100 $Y=577660
X939 1907 2 176 1 INV1S $T=500960 668760 0 0 $X=500960 $Y=668380
X940 1890 2 1898 1 INV1S $T=504060 658680 0 180 $X=502820 $Y=653260
X941 1886 2 1901 1 INV1S $T=505300 638520 0 180 $X=504060 $Y=633100
X942 1914 2 158 1 INV1S $T=504060 709080 1 0 $X=504060 $Y=703660
X943 1885 2 1928 1 INV1S $T=505300 608280 1 0 $X=505300 $Y=602860
X944 1930 2 1915 1 INV1S $T=507160 557880 0 180 $X=505920 $Y=552460
X945 1913 2 181 1 INV1S $T=506540 709080 1 0 $X=506540 $Y=703660
X946 1941 2 1926 1 INV1S $T=510260 567960 1 180 $X=509020 $Y=567580
X947 1944 2 1908 1 INV1S $T=510880 588120 0 180 $X=509640 $Y=582700
X948 1924 2 1937 1 INV1S $T=509640 648600 0 0 $X=509640 $Y=648220
X949 1948 2 178 1 INV1S $T=510880 709080 0 180 $X=509640 $Y=703660
X950 1956 2 1876 1 INV1S $T=511500 628440 0 180 $X=510260 $Y=623020
X951 1920 2 1950 1 INV1S $T=512740 688920 1 180 $X=511500 $Y=688540
X952 1932 2 1960 1 INV1S $T=513360 638520 1 0 $X=513360 $Y=633100
X953 194 2 192 1 INV1S $T=515220 719160 1 0 $X=515220 $Y=713740
X954 1962 2 1918 1 INV1S $T=515840 608280 0 0 $X=515840 $Y=607900
X955 1976 2 1943 1 INV1S $T=518320 557880 1 180 $X=517080 $Y=557500
X956 1977 2 1961 1 INV1S $T=518320 578040 0 180 $X=517080 $Y=572620
X957 1983 2 201 1 INV1S $T=518320 699000 0 0 $X=518320 $Y=698620
X958 1993 2 1935 1 INV1S $T=520800 628440 1 180 $X=519560 $Y=628060
X959 1970 2 1974 1 INV1S $T=520800 588120 1 0 $X=520800 $Y=582700
X960 1995 2 1979 1 INV1S $T=520800 688920 1 0 $X=520800 $Y=683500
X961 2006 2 195 1 INV1S $T=522040 699000 1 180 $X=520800 $Y=698620
X962 2017 2 200 1 INV1S $T=523280 719160 0 180 $X=522040 $Y=713740
X963 2014 2 202 1 INV1S $T=524520 668760 1 180 $X=523280 $Y=668380
X964 2012 2 1972 1 INV1S $T=525140 618360 1 180 $X=523900 $Y=617980
X965 2016 2 1990 1 INV1S $T=525140 648600 1 180 $X=523900 $Y=648220
X966 212 2 1934 1 INV1S $T=526380 608280 0 180 $X=525140 $Y=602860
X967 2018 2 2013 1 INV1S $T=527000 638520 0 180 $X=525760 $Y=633100
X968 2022 2 210 1 INV1S $T=527620 688920 1 180 $X=526380 $Y=688540
X969 2025 2 1987 1 INV1S $T=528240 557880 1 180 $X=527000 $Y=557500
X970 214 2 208 1 INV1S $T=528240 719160 0 180 $X=527000 $Y=713740
X971 2031 2 1978 1 INV1S $T=530100 557880 0 180 $X=528860 $Y=552460
X972 2029 2 1945 1 INV1S $T=530720 678840 1 180 $X=529480 $Y=678460
X973 2026 2 217 1 INV1S $T=529480 719160 1 0 $X=529480 $Y=713740
X974 2044 2 1910 1 INV1S $T=533200 598200 0 180 $X=531960 $Y=592780
X975 2042 2 1997 1 INV1S $T=533200 608280 1 180 $X=531960 $Y=607900
X976 2047 2 1982 1 INV1S $T=533820 638520 0 180 $X=532580 $Y=633100
X977 2035 2 1992 1 INV1S $T=535060 557880 1 180 $X=533820 $Y=557500
X978 2059 2 2000 1 INV1S $T=535680 648600 0 180 $X=534440 $Y=643180
X979 2060 2 1922 1 INV1S $T=536300 618360 1 0 $X=536300 $Y=612940
X980 2083 2 224 1 INV1S $T=537540 688920 0 180 $X=536300 $Y=683500
X981 2072 2 1998 1 INV1S $T=538780 658680 0 180 $X=537540 $Y=653260
X982 2076 2 1939 1 INV1S $T=540640 598200 1 180 $X=539400 $Y=597820
X983 2077 2 223 1 INV1S $T=540640 699000 0 180 $X=539400 $Y=693580
X984 2082 2 2058 1 INV1S $T=541880 598200 1 180 $X=540640 $Y=597820
X985 2074 2 2010 1 INV1S $T=541880 668760 1 180 $X=540640 $Y=668380
X986 2091 2 235 1 INV1S $T=543740 709080 1 180 $X=542500 $Y=708700
X987 2056 2 2068 1 INV1S $T=543740 638520 0 0 $X=543740 $Y=638140
X988 2086 2 2093 1 INV1S $T=543740 688920 1 0 $X=543740 $Y=683500
X989 2099 2 2033 1 INV1S $T=545600 628440 0 180 $X=544360 $Y=623020
X990 239 2 2055 1 INV1S $T=547460 598200 1 180 $X=546220 $Y=597820
X991 2112 2 1949 1 INV1S $T=548080 578040 1 180 $X=546840 $Y=577660
X992 2126 2 2048 1 INV1S $T=549320 658680 0 180 $X=548080 $Y=653260
X993 2105 2 240 1 INV1S $T=549320 688920 1 180 $X=548080 $Y=688540
X994 2102 2 2043 1 INV1S $T=549320 557880 0 0 $X=549320 $Y=557500
X995 2107 2 2036 1 INV1S $T=550560 588120 1 180 $X=549320 $Y=587740
X996 2115 2 2103 1 INV1S $T=551180 678840 0 180 $X=549940 $Y=673420
X997 2122 2 228 1 INV1S $T=552420 709080 0 180 $X=551180 $Y=703660
X998 2118 2 2019 1 INV1S $T=553040 578040 1 180 $X=551800 $Y=577660
X999 2104 2 2080 1 INV1S $T=551800 618360 0 0 $X=551800 $Y=617980
X1000 2114 2 2084 1 INV1S $T=553660 578040 0 180 $X=552420 $Y=572620
X1001 2117 2 2063 1 INV1S $T=554280 668760 0 180 $X=553040 $Y=663340
X1002 2143 2 2111 1 INV1S $T=557380 638520 1 180 $X=556140 $Y=638140
X1003 2140 2 2130 1 INV1S $T=558000 658680 0 180 $X=556760 $Y=653260
X1004 2127 2 2087 1 INV1S $T=557380 719160 1 0 $X=557380 $Y=713740
X1005 2158 2 251 1 INV1S $T=561720 688920 0 0 $X=561720 $Y=688540
X1006 2145 2 2094 1 INV1S $T=562340 567960 0 0 $X=562340 $Y=567580
X1007 2162 2 2095 1 INV1S $T=563580 608280 1 180 $X=562340 $Y=607900
X1008 2167 2 2153 1 INV1S $T=564200 668760 0 180 $X=562960 $Y=663340
X1009 2184 2 2165 1 INV1S $T=566680 628440 1 180 $X=565440 $Y=628060
X1010 2182 2 2132 1 INV1S $T=566680 668760 0 180 $X=565440 $Y=663340
X1011 2178 2 2149 1 INV1S $T=567300 648600 1 180 $X=566060 $Y=648220
X1012 2187 2 2050 1 INV1S $T=567920 588120 0 180 $X=566680 $Y=582700
X1013 2169 2 2124 1 INV1S $T=567920 557880 0 0 $X=567920 $Y=557500
X1014 2195 2 258 1 INV1S $T=569780 688920 1 180 $X=568540 $Y=688540
X1015 2200 2 2159 1 INV1S $T=569780 699000 0 180 $X=568540 $Y=693580
X1016 2196 2 2154 1 INV1S $T=571020 709080 0 180 $X=569780 $Y=703660
X1017 2198 2 2175 1 INV1S $T=572260 658680 0 180 $X=571020 $Y=653260
X1018 2204 2 234 1 INV1S $T=573500 557880 0 180 $X=572260 $Y=552460
X1019 2192 2 2003 1 INV1S $T=572260 578040 0 0 $X=572260 $Y=577660
X1020 2201 2 2032 1 INV1S $T=573500 608280 0 180 $X=572260 $Y=602860
X1021 2202 2 2116 1 INV1S $T=573500 618360 1 180 $X=572260 $Y=617980
X1022 2185 2 1985 1 INV1S $T=574120 598200 1 180 $X=572880 $Y=597820
X1023 2209 2 257 1 INV1S $T=574740 547800 1 0 $X=574740 $Y=542380
X1024 2193 2 2177 1 INV1S $T=574740 628440 1 0 $X=574740 $Y=623020
X1025 2239 2 2212 1 INV1S $T=577220 678840 1 180 $X=575980 $Y=678460
X1026 2210 2 263 1 INV1S $T=575980 709080 0 0 $X=575980 $Y=708700
X1027 2220 2 2194 1 INV1S $T=578460 648600 0 180 $X=577220 $Y=643180
X1028 2217 2 2128 1 INV1S $T=578460 578040 1 0 $X=578460 $Y=572620
X1029 2221 2 2227 1 INV1S $T=583420 658680 0 0 $X=583420 $Y=658300
X1030 239 2 2207 1 INV1S $T=585900 638520 0 180 $X=584660 $Y=633100
X1031 2251 2 2241 1 INV1S $T=586520 699000 0 0 $X=586520 $Y=698620
X1032 2255 2 270 1 INV1S $T=587760 547800 1 0 $X=587760 $Y=542380
X1033 2257 2 268 1 INV1S $T=587760 709080 0 0 $X=587760 $Y=708700
X1034 2259 2 2219 1 INV1S $T=588380 618360 1 0 $X=588380 $Y=612940
X1035 2246 2 2131 1 INV1S $T=589620 608280 0 0 $X=589620 $Y=607900
X1036 2276 2 2188 1 INV1S $T=590860 628440 0 180 $X=589620 $Y=623020
X1037 2271 2 2256 1 INV1S $T=590860 648600 0 0 $X=590860 $Y=648220
X1038 2206 2 2268 1 INV1S $T=590860 668760 1 0 $X=590860 $Y=663340
X1039 2279 2 2250 1 INV1S $T=592100 668760 1 180 $X=590860 $Y=668380
X1040 2272 2 2133 1 INV1S $T=592720 567960 0 180 $X=591480 $Y=562540
X1041 2283 2 2249 1 INV1S $T=592720 578040 1 180 $X=591480 $Y=577660
X1042 2230 2 2247 1 INV1S $T=591480 638520 0 0 $X=591480 $Y=638140
X1043 276 2 274 1 INV1S $T=592720 719160 0 180 $X=591480 $Y=713740
X1044 2297 2 2281 1 INV1S $T=593960 688920 0 180 $X=592720 $Y=683500
X1045 2270 2 231 1 INV1S $T=594580 567960 1 0 $X=594580 $Y=562540
X1046 239 2 2298 1 INV1S $T=595200 588120 0 0 $X=595200 $Y=587740
X1047 2304 2 2309 1 INV1S $T=598300 678840 1 0 $X=598300 $Y=673420
X1048 2321 2 2197 1 INV1S $T=600160 608280 0 180 $X=598920 $Y=602860
X1049 2315 2 2253 1 INV1S $T=600160 628440 0 180 $X=598920 $Y=623020
X1050 2285 2 2295 1 INV1S $T=598920 638520 0 0 $X=598920 $Y=638140
X1051 2336 2 2300 1 INV1S $T=603260 678840 0 180 $X=602020 $Y=673420
X1052 2264 2 2311 1 INV1S $T=602020 699000 1 0 $X=602020 $Y=693580
X1053 2327 2 2073 1 INV1S $T=603880 557880 0 180 $X=602640 $Y=552460
X1054 2332 2 2173 1 INV1S $T=603880 588120 1 180 $X=602640 $Y=587740
X1055 2324 2 2280 1 INV1S $T=603880 709080 0 180 $X=602640 $Y=703660
X1056 2326 2 279 1 INV1S $T=605120 547800 1 180 $X=603880 $Y=547420
X1057 2318 2 2267 1 INV1S $T=604500 658680 1 0 $X=604500 $Y=653260
X1058 2317 2 2340 1 INV1S $T=605740 638520 1 0 $X=605740 $Y=633100
X1059 2325 2 2334 1 INV1S $T=606980 658680 1 0 $X=606980 $Y=653260
X1060 2346 2 2288 1 INV1S $T=607600 678840 0 0 $X=607600 $Y=678460
X1061 2358 2 2299 1 INV1S $T=609460 668760 1 0 $X=609460 $Y=663340
X1062 2341 2 2328 1 INV1S $T=610700 628440 1 0 $X=610700 $Y=623020
X1063 2362 2 2141 1 INV1S $T=612560 608280 0 180 $X=611320 $Y=602860
X1064 2352 2 2354 1 INV1S $T=611320 688920 1 0 $X=611320 $Y=683500
X1065 2371 2 2342 1 INV1S $T=612560 699000 1 180 $X=611320 $Y=698620
X1066 2366 2 2350 1 INV1S $T=612560 618360 1 0 $X=612560 $Y=612940
X1067 2368 2 2218 1 INV1S $T=613180 567960 1 0 $X=613180 $Y=562540
X1068 2381 2 267 1 INV1S $T=615660 547800 0 0 $X=615660 $Y=547420
X1069 2344 2 2260 1 INV1S $T=616280 567960 0 0 $X=616280 $Y=567580
X1070 2389 2 288 1 INV1S $T=619380 547800 1 180 $X=618140 $Y=547420
X1071 2082 2 2379 1 INV1S $T=618140 658680 1 0 $X=618140 $Y=653260
X1072 2363 2 2236 1 INV1S $T=620000 578040 1 0 $X=620000 $Y=572620
X1073 2382 2 2378 1 INV1S $T=621240 668760 0 0 $X=621240 $Y=668380
X1074 2417 2 2399 1 INV1S $T=622480 699000 0 0 $X=622480 $Y=698620
X1075 2416 2 2430 1 INV1S $T=624960 588120 0 0 $X=624960 $Y=587740
X1076 2420 2 2373 1 INV1S $T=624960 688920 0 0 $X=624960 $Y=688540
X1077 2423 2 2409 1 INV1S $T=626200 699000 1 180 $X=624960 $Y=698620
X1078 2428 2 2349 1 INV1S $T=626820 628440 0 180 $X=625580 $Y=623020
X1079 2429 2 2412 1 INV1S $T=626820 638520 0 180 $X=625580 $Y=633100
X1080 2375 2 2434 1 INV1S $T=626820 578040 1 0 $X=626820 $Y=572620
X1081 2375 2 2435 1 INV1S $T=626820 608280 1 0 $X=626820 $Y=602860
X1082 2439 2 2415 1 INV1S $T=628060 719160 0 180 $X=626820 $Y=713740
X1083 2433 2 2277 1 INV1S $T=627440 567960 1 0 $X=627440 $Y=562540
X1084 2440 2 2331 1 INV1S $T=628680 588120 1 180 $X=627440 $Y=587740
X1085 2442 2 2357 1 INV1S $T=629300 678840 0 180 $X=628060 $Y=673420
X1086 2425 2 2443 1 INV1S $T=628680 688920 0 0 $X=628680 $Y=688540
X1087 2441 2 2411 1 INV1S $T=629300 608280 1 0 $X=629300 $Y=602860
X1088 2436 2 2390 1 INV1S $T=630540 608280 1 180 $X=629300 $Y=607900
X1089 2458 2 2191 1 INV1S $T=633020 557880 0 180 $X=631780 $Y=552460
X1090 2465 2 2438 1 INV1S $T=634260 638520 0 180 $X=633020 $Y=633100
X1091 2466 2 2403 1 INV1S $T=635500 648600 1 180 $X=634260 $Y=648220
X1092 2463 2 2427 1 INV1S $T=634260 658680 0 0 $X=634260 $Y=658300
X1093 311 2 307 1 INV1S $T=636120 719160 0 180 $X=634880 $Y=713740
X1094 2447 2 2248 1 INV1S $T=637980 547800 1 180 $X=636740 $Y=547420
X1095 2469 2 2474 1 INV1S $T=637980 648600 1 180 $X=636740 $Y=648220
X1096 2449 2 2476 1 INV1S $T=637980 668760 0 0 $X=637980 $Y=668380
X1097 2486 2 2303 1 INV1S $T=640460 567960 0 0 $X=640460 $Y=567580
X1098 2504 2 2432 1 INV1S $T=643560 598200 0 180 $X=642320 $Y=592780
X1099 2490 2 2464 1 INV1S $T=643560 678840 1 180 $X=642320 $Y=678460
X1100 2499 2 2477 1 INV1S $T=643560 699000 0 180 $X=642320 $Y=693580
X1101 2508 2 314 1 INV1S $T=644180 709080 1 180 $X=642940 $Y=708700
X1102 2506 2 2485 1 INV1S $T=645420 588120 0 0 $X=645420 $Y=587740
X1103 2513 2 2355 1 INV1S $T=646660 608280 0 180 $X=645420 $Y=602860
X1104 2518 2 2384 1 INV1S $T=647280 709080 1 180 $X=646040 $Y=708700
X1105 317 2 2516 1 INV1S $T=646660 547800 0 0 $X=646660 $Y=547420
X1106 2517 2 2503 1 INV1S $T=647900 648600 0 180 $X=646660 $Y=643180
X1107 2519 2 315 1 INV1S $T=649140 578040 1 180 $X=647900 $Y=577660
X1108 2545 2 2511 1 INV1S $T=649760 678840 1 180 $X=648520 $Y=678460
X1109 2521 2 2408 1 INV1S $T=650380 618360 1 180 $X=649140 $Y=617980
X1110 2523 2 2396 1 INV1S $T=651000 608280 1 180 $X=649760 $Y=607900
X1111 2533 2 2522 1 INV1S $T=651620 688920 0 180 $X=650380 $Y=683500
X1112 2529 2 2501 1 INV1S $T=652240 588120 1 180 $X=651000 $Y=587740
X1113 2531 2 2502 1 INV1S $T=652240 668760 0 180 $X=651000 $Y=663340
X1114 2538 2 319 1 INV1S $T=652240 709080 1 180 $X=651000 $Y=708700
X1115 2532 2 2530 1 INV1S $T=651620 709080 1 0 $X=651620 $Y=703660
X1116 2536 2 2535 1 INV1S $T=653480 638520 0 0 $X=653480 $Y=638140
X1117 2554 2 2534 1 INV1S $T=655340 588120 0 180 $X=654100 $Y=582700
X1118 2553 2 320 1 INV1S $T=656580 567960 1 180 $X=655340 $Y=567580
X1119 2566 2 328 1 INV1S $T=658440 567960 0 180 $X=657200 $Y=562540
X1120 2563 2 2473 1 INV1S $T=658440 628440 1 180 $X=657200 $Y=628060
X1121 332 2 2542 1 INV1S $T=659060 547800 0 180 $X=657820 $Y=542380
X1122 2569 2 2356 1 INV1S $T=659680 618360 0 180 $X=658440 $Y=612940
X1123 2562 2 2487 1 INV1S $T=659680 699000 1 180 $X=658440 $Y=698620
X1124 2581 2 2543 1 INV1S $T=660300 688920 0 180 $X=659060 $Y=683500
X1125 2573 2 333 1 INV1S $T=660300 709080 1 180 $X=659060 $Y=708700
X1126 2576 2 2540 1 INV1S $T=662160 658680 1 180 $X=660920 $Y=658300
X1127 2571 2 334 1 INV1S $T=665260 578040 0 180 $X=664020 $Y=572620
X1128 336 2 2575 1 INV1S $T=665880 557880 0 0 $X=665880 $Y=557500
X1129 2515 2 2588 1 INV1S $T=667120 598200 1 180 $X=665880 $Y=597820
X1130 2598 2 2478 1 INV1S $T=668360 628440 0 180 $X=667120 $Y=623020
X1131 2593 2 2551 1 INV1S $T=668980 688920 1 180 $X=667740 $Y=688540
X1132 2596 2 2498 1 INV1S $T=669600 638520 0 180 $X=668360 $Y=633100
X1133 2594 2 2539 1 INV1S $T=671460 567960 1 180 $X=670220 $Y=567580
X1134 2599 2 2597 1 INV1S $T=671460 588120 0 180 $X=670220 $Y=582700
X1135 2603 2 2577 1 INV1S $T=672080 658680 0 180 $X=670840 $Y=653260
X1136 2609 2 2570 1 INV1S $T=674560 688920 1 180 $X=673320 $Y=688540
X1137 2612 2 2595 1 INV1S $T=675800 709080 0 180 $X=674560 $Y=703660
X1138 343 2 2605 1 INV1S $T=675800 547800 0 0 $X=675800 $Y=547420
X1139 344 2 2617 1 INV1S $T=677040 547800 0 0 $X=677040 $Y=547420
X1140 2620 2 2568 1 INV1S $T=678280 668760 0 180 $X=677040 $Y=663340
X1141 2602 2 346 1 INV1S $T=677660 567960 1 0 $X=677660 $Y=562540
X1142 353 2 2583 1 INV1S $T=686960 557880 0 180 $X=685720 $Y=552460
X1143 2645 2 2640 1 INV1S $T=686960 598200 0 180 $X=685720 $Y=592780
X1144 2661 2 352 1 INV1S $T=687580 709080 1 180 $X=686340 $Y=708700
X1145 2646 2 354 1 INV1S $T=688820 678840 0 0 $X=688820 $Y=678460
X1146 2652 2 355 1 INV1S $T=688820 688920 0 0 $X=688820 $Y=688540
X1147 2670 2 2672 1 INV1S $T=692540 567960 0 180 $X=691300 $Y=562540
X1148 2680 2 2665 1 INV1S $T=693160 578040 1 0 $X=693160 $Y=572620
X1149 2691 2 2666 1 INV1S $T=695020 557880 0 180 $X=693780 $Y=552460
X1150 2686 2 2674 1 INV1S $T=696260 557880 1 180 $X=695020 $Y=557500
X1151 2698 2 2676 1 INV1S $T=696260 578040 0 180 $X=695020 $Y=572620
X1152 2660 2 350 1 INV1S $T=695020 699000 1 0 $X=695020 $Y=693580
X1153 2656 2 2688 1 INV1S $T=696880 618360 0 180 $X=695640 $Y=612940
X1154 2642 2 2687 1 INV1S $T=697500 628440 0 0 $X=697500 $Y=628060
X1155 2655 2 2705 1 INV1S $T=698120 557880 0 0 $X=698120 $Y=557500
X1156 2629 2 2703 1 INV1S $T=698120 598200 0 0 $X=698120 $Y=597820
X1157 2662 2 2745 1 INV1S $T=702460 628440 1 0 $X=702460 $Y=623020
X1158 371 2 2731 1 INV1S $T=703700 709080 1 180 $X=702460 $Y=708700
X1159 2752 2 2730 1 INV1S $T=704940 547800 1 180 $X=703700 $Y=547420
X1160 2647 2 2743 1 INV1S $T=704940 578040 1 180 $X=703700 $Y=577660
X1161 2761 2 2748 1 INV1S $T=707420 588120 0 180 $X=706180 $Y=582700
X1162 2727 2 2755 1 INV1S $T=707420 638520 0 180 $X=706180 $Y=633100
X1163 2759 2 2721 1 INV1S $T=707420 688920 0 180 $X=706180 $Y=683500
X1164 2704 2 2777 1 INV1S $T=706800 608280 0 0 $X=706800 $Y=607900
X1165 2758 2 2766 1 INV1S $T=706800 628440 0 0 $X=706800 $Y=628060
X1166 2767 2 2775 1 INV1S $T=707420 709080 1 0 $X=707420 $Y=703660
X1167 2719 2 2778 1 INV1S $T=708660 638520 0 0 $X=708660 $Y=638140
X1168 2770 2 2780 1 INV1S $T=708660 699000 1 0 $X=708660 $Y=693580
X1169 2702 2 2786 1 INV1S $T=709900 567960 0 0 $X=709900 $Y=567580
X1170 2772 2 2809 1 INV1S $T=711140 628440 1 0 $X=711140 $Y=623020
X1171 2656 2 2805 1 INV1S $T=711760 618360 1 0 $X=711760 $Y=612940
X1172 2806 2 2791 1 INV1S $T=713620 648600 1 180 $X=712380 $Y=648220
X1173 2774 2 2821 1 INV1S $T=714240 598200 0 0 $X=714240 $Y=597820
X1174 2766 2 2826 1 INV1S $T=714240 638520 1 0 $X=714240 $Y=633100
X1175 2824 2 2776 1 INV1S $T=715480 688920 0 180 $X=714240 $Y=683500
X1176 2824 2 2789 1 INV1S $T=716100 699000 1 180 $X=714860 $Y=698620
X1177 2824 2 2796 1 INV1S $T=716720 709080 0 180 $X=715480 $Y=703660
X1178 2842 2 2852 1 INV1S $T=717960 578040 1 0 $X=717960 $Y=572620
X1179 2828 2 2863 1 INV1S $T=719820 668760 1 0 $X=719820 $Y=663340
X1180 2856 2 2879 1 INV1S $T=721060 658680 1 0 $X=721060 $Y=653260
X1181 2861 2 2868 1 INV1S $T=721680 567960 0 0 $X=721680 $Y=567580
X1182 2823 2 2892 1 INV1S $T=721680 668760 1 0 $X=721680 $Y=663340
X1183 2637 2 2893 1 INV1S $T=722300 578040 0 0 $X=722300 $Y=577660
X1184 2858 2 2885 1 INV1S $T=722920 688920 0 0 $X=722920 $Y=688540
X1185 366 2 2915 1 INV1S $T=722920 709080 0 0 $X=722920 $Y=708700
X1186 2855 2 2877 1 INV1S $T=723540 567960 0 0 $X=723540 $Y=567580
X1187 2893 2 2906 1 INV1S $T=724780 578040 0 0 $X=724780 $Y=577660
X1188 2899 2 2907 1 INV1S $T=724780 678840 0 0 $X=724780 $Y=678460
X1189 2736 2 2735 1 INV1S $T=726020 578040 1 0 $X=726020 $Y=572620
X1190 2866 2 2929 1 INV1S $T=726640 608280 1 0 $X=726640 $Y=602860
X1191 2893 2 2925 1 INV1S $T=727260 588120 1 0 $X=727260 $Y=582700
X1192 2925 2 2825 1 INV1S $T=728500 588120 1 180 $X=727260 $Y=587740
X1193 2929 2 2850 1 INV1S $T=728500 598200 1 180 $X=727260 $Y=597820
X1194 396 2 2920 1 INV1S $T=728500 678840 1 180 $X=727260 $Y=678460
X1195 2922 2 2883 1 INV1S $T=730360 578040 0 180 $X=729120 $Y=572620
X1196 2930 2 2945 1 INV1S $T=729740 678840 0 0 $X=729740 $Y=678460
X1197 2916 2 2941 1 INV1S $T=730360 547800 0 0 $X=730360 $Y=547420
X1198 2960 2 2811 1 INV1S $T=732220 598200 1 180 $X=730980 $Y=597820
X1199 2951 2 2946 1 INV1S $T=732220 658680 1 180 $X=730980 $Y=658300
X1200 2842 2 2957 1 INV1S $T=731600 588120 1 0 $X=731600 $Y=582700
X1201 2870 2 2940 1 INV1S $T=732840 598200 0 180 $X=731600 $Y=592780
X1202 2924 2 2950 1 INV1S $T=732840 547800 0 0 $X=732840 $Y=547420
X1203 2952 2 2939 1 INV1S $T=733460 668760 1 0 $X=733460 $Y=663340
X1204 401 2 3002 1 INV1S $T=735320 709080 0 0 $X=735320 $Y=708700
X1205 2968 2 2995 1 INV1S $T=735940 678840 0 0 $X=735940 $Y=678460
X1206 2808 2 2982 1 INV1S $T=737180 567960 1 0 $X=737180 $Y=562540
X1207 2999 2 3004 1 INV1S $T=738420 618360 0 0 $X=738420 $Y=617980
X1208 2979 2 2996 1 INV1S $T=738420 709080 1 0 $X=738420 $Y=703660
X1209 2976 2 3006 1 INV1S $T=739040 598200 1 0 $X=739040 $Y=592780
X1210 2890 2 3023 1 INV1S $T=741520 547800 0 0 $X=741520 $Y=547420
X1211 384 2 2973 1 INV1S $T=742760 678840 0 180 $X=741520 $Y=673420
X1212 2992 2 3029 1 INV1S $T=741520 699000 1 0 $X=741520 $Y=693580
X1213 3015 2 3026 1 INV1S $T=742140 598200 0 0 $X=742140 $Y=597820
X1214 3027 2 3017 1 INV1S $T=743380 688920 0 180 $X=742140 $Y=683500
X1215 3003 2 3049 1 INV1S $T=742760 547800 0 0 $X=742760 $Y=547420
X1216 2991 2 3033 1 INV1S $T=742760 678840 0 0 $X=742760 $Y=678460
X1217 3012 2 3046 1 INV1S $T=743380 628440 0 0 $X=743380 $Y=628060
X1218 2988 2 3021 1 INV1S $T=745860 658680 0 180 $X=744620 $Y=653260
X1219 2844 2 3051 1 INV1S $T=745860 567960 1 0 $X=745860 $Y=562540
X1220 3040 2 3059 1 INV1S $T=745860 598200 1 0 $X=745860 $Y=592780
X1221 2913 2 3053 1 INV1S $T=747720 658680 1 180 $X=746480 $Y=658300
X1222 3057 2 3044 1 INV1S $T=747720 709080 1 180 $X=746480 $Y=708700
X1223 3063 2 3050 1 INV1S $T=747720 557880 0 0 $X=747720 $Y=557500
X1224 3042 2 3070 1 INV1S $T=748340 628440 1 0 $X=748340 $Y=623020
X1225 3043 2 3081 1 INV1S $T=749580 688920 0 0 $X=749580 $Y=688540
X1226 3072 2 3095 1 INV1S $T=750820 699000 1 0 $X=750820 $Y=693580
X1227 3079 2 3090 1 INV1S $T=751440 648600 0 0 $X=751440 $Y=648220
X1228 3048 2 3061 1 INV1S $T=752680 658680 0 180 $X=751440 $Y=653260
X1229 3097 2 3069 1 INV1S $T=753300 598200 1 0 $X=753300 $Y=592780
X1230 2975 2 3117 1 INV1S $T=753920 578040 1 0 $X=753920 $Y=572620
X1231 422 2 2994 1 INV1S $T=755780 719160 0 180 $X=754540 $Y=713740
X1232 3039 2 3113 1 INV1S $T=756400 699000 0 0 $X=756400 $Y=698620
X1233 3120 2 3109 1 INV1S $T=758260 608280 1 180 $X=757020 $Y=607900
X1234 3102 2 3127 1 INV1S $T=757640 628440 1 0 $X=757640 $Y=623020
X1235 422 2 3132 1 INV1S $T=758260 719160 1 0 $X=758260 $Y=713740
X1236 417 2 3143 1 INV1S $T=759500 719160 1 0 $X=759500 $Y=713740
X1237 3115 2 3130 1 INV1S $T=762600 618360 0 180 $X=761360 $Y=612940
X1238 3058 2 3151 1 INV1S $T=761980 588120 1 0 $X=761980 $Y=582700
X1239 3136 2 3159 1 INV1S $T=763220 628440 1 0 $X=763220 $Y=623020
X1240 2671 2 3162 1 INV1S $T=763840 588120 1 0 $X=763840 $Y=582700
X1241 2785 2 3166 1 INV1S $T=764460 628440 1 0 $X=764460 $Y=623020
X1242 3158 2 3175 1 INV1S $T=765700 658680 1 0 $X=765700 $Y=653260
X1243 3171 2 3177 1 INV1S $T=766320 608280 0 0 $X=766320 $Y=607900
X1244 2802 2 3188 1 INV1S $T=768800 699000 1 180 $X=767560 $Y=698620
X1245 3141 2 3192 1 INV1S $T=767560 709080 1 0 $X=767560 $Y=703660
X1246 2839 2 3205 1 INV1S $T=768800 678840 0 0 $X=768800 $Y=678460
X1247 3129 2 3197 1 INV1S $T=771900 578040 1 180 $X=770660 $Y=577660
X1248 2822 2 3226 1 INV1S $T=770660 628440 1 0 $X=770660 $Y=623020
X1249 3193 2 3216 1 INV1S $T=771280 588120 0 0 $X=771280 $Y=587740
X1250 3052 2 3223 1 INV1S $T=771900 567960 0 0 $X=771900 $Y=567580
X1251 2886 2 3230 1 INV1S $T=772520 608280 0 0 $X=772520 $Y=607900
X1252 3152 2 3228 1 INV1S $T=772520 648600 1 0 $X=772520 $Y=643180
X1253 3172 2 3225 1 INV1S $T=774380 709080 0 180 $X=773140 $Y=703660
X1254 3220 2 3237 1 INV1S $T=773760 709080 0 0 $X=773760 $Y=708700
X1255 3206 2 3238 1 INV1S $T=773760 719160 1 0 $X=773760 $Y=713740
X1256 3207 2 3249 1 INV1S $T=775000 567960 1 0 $X=775000 $Y=562540
X1257 3134 2 3234 1 INV1S $T=776860 588120 1 0 $X=776860 $Y=582700
X1258 3239 2 3268 1 INV1S $T=777480 567960 1 0 $X=777480 $Y=562540
X1259 3160 2 3260 1 INV1S $T=777480 608280 1 0 $X=777480 $Y=602860
X1260 3180 2 3264 1 INV1S $T=778100 648600 1 0 $X=778100 $Y=643180
X1261 3088 2 3267 1 INV1S $T=778720 688920 1 0 $X=778720 $Y=683500
X1262 3251 2 3273 1 INV1S $T=779340 628440 1 0 $X=779340 $Y=623020
X1263 3219 2 3274 1 INV1S $T=779960 688920 1 0 $X=779960 $Y=683500
X1264 433 2 432 1 INV1S $T=781200 719160 0 180 $X=779960 $Y=713740
X1265 3291 2 3296 1 INV1S $T=783060 678840 0 0 $X=783060 $Y=678460
X1266 2840 2 3285 1 INV1S $T=784300 709080 1 180 $X=783060 $Y=708700
X1267 3304 2 3311 1 INV1S $T=786160 578040 1 0 $X=786160 $Y=572620
X1268 3320 2 3341 1 INV1S $T=789880 628440 0 0 $X=789880 $Y=628060
X1269 437 2 3328 1 INV1S $T=790500 547800 1 0 $X=790500 $Y=542380
X1270 3312 2 3346 1 INV1S $T=790500 588120 1 0 $X=790500 $Y=582700
X1271 3091 2 3350 1 INV1S $T=791740 638520 1 0 $X=791740 $Y=633100
X1272 3266 2 3372 1 INV1S $T=792980 638520 1 0 $X=792980 $Y=633100
X1273 3352 2 3358 1 INV1S $T=792980 699000 0 0 $X=792980 $Y=698620
X1274 3259 2 3353 1 INV1S $T=792980 719160 1 0 $X=792980 $Y=713740
X1275 3292 2 3364 1 INV1S $T=793600 688920 1 0 $X=793600 $Y=683500
X1276 3298 2 3355 1 INV1S $T=794220 588120 0 0 $X=794220 $Y=587740
X1277 3242 2 3384 1 INV1S $T=794840 688920 1 0 $X=794840 $Y=683500
X1278 3339 2 3381 1 INV1S $T=795460 557880 1 0 $X=795460 $Y=552460
X1279 3001 2 3344 1 INV1S $T=795460 709080 0 0 $X=795460 $Y=708700
X1280 3382 2 3377 1 INV1S $T=796700 578040 0 0 $X=796700 $Y=577660
X1281 3365 2 3367 1 INV1S $T=800420 557880 1 180 $X=799180 $Y=557500
X1282 3404 2 3397 1 INV1S $T=801040 578040 1 180 $X=799800 $Y=577660
X1283 3314 2 3398 1 INV1S $T=802900 557880 1 0 $X=802900 $Y=552460
X1284 3343 2 3440 1 INV1S $T=803520 638520 0 0 $X=803520 $Y=638140
X1285 3279 2 3456 1 INV1S $T=804140 648600 0 0 $X=804140 $Y=648220
X1286 3431 2 3443 1 INV1S $T=805380 608280 0 0 $X=805380 $Y=607900
X1287 3447 2 3458 1 INV1S $T=806620 567960 0 0 $X=806620 $Y=567580
X1288 3453 2 3396 1 INV1S $T=807860 608280 1 0 $X=807860 $Y=602860
X1289 3217 2 3463 1 INV1S $T=807860 648600 1 0 $X=807860 $Y=643180
X1290 3468 2 3457 1 INV1S $T=809720 688920 0 180 $X=808480 $Y=683500
X1291 3415 2 3459 1 INV1S $T=811580 618360 0 180 $X=810340 $Y=612940
X1292 3437 2 3475 1 INV1S $T=810960 678840 1 0 $X=810960 $Y=673420
X1293 3370 2 3481 1 INV1S $T=811580 648600 0 0 $X=811580 $Y=648220
X1294 3469 2 3487 1 INV1S $T=812200 618360 0 0 $X=812200 $Y=617980
X1295 3449 2 3490 1 INV1S $T=812820 618360 1 0 $X=812820 $Y=612940
X1296 3442 2 3489 1 INV1S $T=812820 678840 0 0 $X=812820 $Y=678460
X1297 3485 2 3497 1 INV1S $T=814060 699000 1 0 $X=814060 $Y=693580
X1298 3401 2 3508 1 INV1S $T=814680 668760 0 0 $X=814680 $Y=668380
X1299 3424 2 3486 1 INV1S $T=815300 567960 0 0 $X=815300 $Y=567580
X1300 3418 2 3501 1 INV1S $T=815300 638520 1 0 $X=815300 $Y=633100
X1301 3451 2 3520 1 INV1S $T=817780 658680 0 0 $X=817780 $Y=658300
X1302 3488 2 3525 1 INV1S $T=818400 709080 1 0 $X=818400 $Y=703660
X1303 3522 2 3528 1 INV1S $T=820880 618360 1 0 $X=820880 $Y=612940
X1304 3464 2 3537 1 INV1S $T=823360 709080 1 0 $X=823360 $Y=703660
X1305 3517 2 3551 1 INV1S $T=825840 699000 0 0 $X=825840 $Y=698620
X1306 3542 2 3564 1 INV1S $T=830800 618360 0 0 $X=830800 $Y=617980
X1307 3582 2 3576 1 INV1S $T=834520 688920 1 180 $X=833280 $Y=688540
X1308 3571 2 3587 1 INV1S $T=834520 618360 1 0 $X=834520 $Y=612940
X1309 3597 2 3593 1 INV1S $T=838860 688920 1 180 $X=837620 $Y=688540
X1310 479 2 3591 1 INV1S $T=838860 688920 1 0 $X=838860 $Y=683500
X1311 3609 2 3610 1 INV1S $T=839480 608280 1 0 $X=839480 $Y=602860
X1312 3596 2 3608 1 INV1S $T=840720 699000 1 180 $X=839480 $Y=698620
X1313 3589 2 3614 1 INV1S $T=840100 588120 0 0 $X=840100 $Y=587740
X1314 3605 2 3643 1 INV1S $T=840720 688920 1 0 $X=840720 $Y=683500
X1315 3628 2 3606 1 INV1S $T=842580 618360 1 180 $X=841340 $Y=617980
X1316 3626 2 3631 1 INV1S $T=842580 557880 0 0 $X=842580 $Y=557500
X1317 3622 2 3632 1 INV1S $T=842580 678840 1 0 $X=842580 $Y=673420
X1318 3621 2 3661 1 INV1S $T=846300 598200 0 0 $X=846300 $Y=597820
X1319 3633 2 3665 1 INV1S $T=847540 578040 1 0 $X=847540 $Y=572620
X1320 3650 2 3649 1 INV1S $T=847540 668760 0 0 $X=847540 $Y=668380
X1321 3645 2 3668 1 INV1S $T=848160 567960 1 0 $X=848160 $Y=562540
X1322 3669 2 3677 1 INV1S $T=848780 578040 1 0 $X=848780 $Y=572620
X1323 3635 2 3679 1 INV1S $T=850020 699000 1 0 $X=850020 $Y=693580
X1324 3659 2 3666 1 INV1S $T=850640 598200 1 0 $X=850640 $Y=592780
X1325 3667 2 3691 1 INV1S $T=852500 547800 1 0 $X=852500 $Y=542380
X1326 3651 2 3693 1 INV1S $T=853120 567960 0 0 $X=853120 $Y=567580
X1327 3653 2 3686 1 INV1S $T=856220 557880 1 180 $X=854980 $Y=557500
X1328 505 2 509 1 INV1S $T=864280 547800 0 0 $X=864280 $Y=547420
X1329 3730 2 3736 1 INV1S $T=866760 547800 0 0 $X=866760 $Y=547420
X1330 510 2 3715 1 INV1S $T=868000 719160 0 180 $X=866760 $Y=713740
X1331 3731 2 3732 1 INV1S $T=868620 638520 0 180 $X=867380 $Y=633100
X1332 514 2 3723 1 INV1S $T=870480 719160 0 180 $X=869240 $Y=713740
X1333 3746 2 3754 1 INV1S $T=871100 648600 0 180 $X=869860 $Y=643180
X1334 3762 2 3755 1 INV1S $T=871100 658680 0 180 $X=869860 $Y=653260
X1335 3751 2 3777 1 INV1S $T=871100 557880 0 0 $X=871100 $Y=557500
X1336 3773 2 3770 1 INV1S $T=873580 648600 1 180 $X=872340 $Y=648220
X1337 3771 2 3767 1 INV1S $T=874820 709080 0 180 $X=873580 $Y=703660
X1338 3776 2 3782 1 INV1S $T=874200 557880 1 0 $X=874200 $Y=552460
X1339 3768 2 3801 1 INV1S $T=876060 557880 0 0 $X=876060 $Y=557500
X1340 3817 2 3781 1 INV1S $T=878540 658680 1 180 $X=877300 $Y=658300
X1341 3788 2 3800 1 INV1S $T=877300 719160 1 0 $X=877300 $Y=713740
X1342 3794 2 3797 1 INV1S $T=879160 658680 0 180 $X=877920 $Y=653260
X1343 3663 2 3757 1 INV1S $T=879780 648600 0 180 $X=878540 $Y=643180
X1344 522 2 3820 1 INV1S $T=879160 709080 0 0 $X=879160 $Y=708700
X1345 3833 2 3838 1 INV1S $T=883500 638520 0 0 $X=883500 $Y=638140
X1346 3819 2 3845 1 INV1S $T=884120 658680 1 0 $X=884120 $Y=653260
X1347 3832 2 3875 1 INV1S $T=887220 588120 1 0 $X=887220 $Y=582700
X1348 3784 2 3863 1 INV1S $T=887840 557880 0 0 $X=887840 $Y=557500
X1349 3828 2 3858 1 INV1S $T=890940 638520 1 180 $X=889700 $Y=638140
X1350 3884 2 3837 1 INV1S $T=890940 658680 0 180 $X=889700 $Y=653260
X1351 3877 2 3894 1 INV1S $T=890940 557880 0 0 $X=890940 $Y=557500
X1352 3809 2 3852 1 INV1S $T=890940 648600 1 0 $X=890940 $Y=643180
X1353 3836 2 3883 1 INV1S $T=893420 567960 1 180 $X=892180 $Y=567580
X1354 3892 2 3857 1 INV1S $T=894040 688920 1 180 $X=892800 $Y=688540
X1355 3898 2 3881 1 INV1S $T=894660 688920 0 180 $X=893420 $Y=683500
X1356 3796 2 3922 1 INV1S $T=896520 578040 0 0 $X=896520 $Y=577660
X1357 3910 2 3915 1 INV1S $T=897760 658680 1 180 $X=896520 $Y=658300
X1358 3906 2 3935 1 INV1S $T=897140 567960 0 0 $X=897140 $Y=567580
X1359 3885 2 3939 1 INV1S $T=899000 638520 0 0 $X=899000 $Y=638140
X1360 3909 2 3958 1 INV1S $T=899000 648600 1 0 $X=899000 $Y=643180
X1361 3867 2 3943 1 INV1S $T=899620 567960 0 0 $X=899620 $Y=567580
X1362 3944 2 3927 1 INV1S $T=900860 688920 1 180 $X=899620 $Y=688540
X1363 547 2 3926 1 INV1S $T=902720 547800 1 180 $X=901480 $Y=547420
X1364 3956 2 3950 1 INV1S $T=902720 588120 0 180 $X=901480 $Y=582700
X1365 3889 2 3974 1 INV1S $T=902100 598200 1 0 $X=902100 $Y=592780
X1366 3822 2 3946 1 INV1S $T=902720 578040 0 0 $X=902720 $Y=577660
X1367 3952 2 3959 1 INV1S $T=903340 638520 0 0 $X=903340 $Y=638140
X1368 3963 2 3984 1 INV1S $T=905200 709080 1 0 $X=905200 $Y=703660
X1369 3972 2 3985 1 INV1S $T=905820 567960 0 0 $X=905820 $Y=567580
X1370 549 2 3980 1 INV1S $T=905820 699000 0 0 $X=905820 $Y=698620
X1371 3981 2 3973 1 INV1S $T=908300 588120 0 180 $X=907060 $Y=582700
X1372 3999 2 3998 1 INV1S $T=910780 567960 1 180 $X=909540 $Y=567580
X1373 4009 2 4001 1 INV1S $T=911400 638520 1 180 $X=910160 $Y=638140
X1374 3975 2 4002 1 INV1S $T=911400 648600 1 180 $X=910160 $Y=648220
X1375 4018 2 3976 1 INV1S $T=912640 638520 1 180 $X=911400 $Y=638140
X1376 555 2 564 1 INV1S $T=912020 547800 1 0 $X=912020 $Y=542380
X1377 4007 2 4005 1 INV1S $T=912020 588120 0 0 $X=912020 $Y=587740
X1378 4048 2 562 1 INV1S $T=915740 598200 1 180 $X=914500 $Y=597820
X1379 4028 2 4012 1 INV1S $T=915120 567960 1 0 $X=915120 $Y=562540
X1380 4042 2 4034 1 INV1S $T=916980 688920 0 180 $X=915740 $Y=683500
X1381 4046 2 4049 1 INV1S $T=916980 567960 1 0 $X=916980 $Y=562540
X1382 4044 2 4055 1 INV1S $T=917600 648600 1 0 $X=917600 $Y=643180
X1383 4064 2 4072 1 INV1S $T=920080 648600 1 0 $X=920080 $Y=643180
X1384 566 2 4066 1 INV1S $T=921320 699000 1 180 $X=920080 $Y=698620
X1385 4083 2 4071 1 INV1S $T=921940 628440 1 180 $X=920700 $Y=628060
X1386 3908 2 4103 1 INV1S $T=923800 567960 0 0 $X=923800 $Y=567580
X1387 4030 2 4094 1 INV1S $T=925660 678840 1 180 $X=924420 $Y=678460
X1388 4051 2 4109 1 INV1S $T=925660 709080 1 0 $X=925660 $Y=703660
X1389 3901 2 4116 1 INV1S $T=926280 567960 0 0 $X=926280 $Y=567580
X1390 4108 2 4114 1 INV1S $T=928140 588120 0 180 $X=926900 $Y=582700
X1391 4124 2 4115 1 INV1S $T=928760 628440 1 180 $X=927520 $Y=628060
X1392 4076 2 4097 1 INV1S $T=929380 588120 0 180 $X=928140 $Y=582700
X1393 4130 2 4137 1 INV1S $T=929380 547800 0 0 $X=929380 $Y=547420
X1394 4135 2 4134 1 INV1S $T=930620 628440 1 180 $X=929380 $Y=628060
X1395 4127 2 4153 1 INV1S $T=931240 588120 0 0 $X=931240 $Y=587740
X1396 4118 2 4132 1 INV1S $T=932480 638520 0 180 $X=931240 $Y=633100
X1397 4119 2 4120 1 INV1S $T=932480 557880 0 0 $X=932480 $Y=557500
X1398 4105 2 4155 1 INV1S $T=936200 557880 1 180 $X=934960 $Y=557500
X1399 4165 2 4150 1 INV1S $T=939300 638520 0 180 $X=938060 $Y=633100
X1400 4174 2 4160 1 INV1S $T=939920 628440 0 0 $X=939920 $Y=628060
X1401 4190 2 4180 1 INV1S $T=942400 699000 0 180 $X=941160 $Y=693580
X1402 4177 2 4187 1 INV1S $T=941780 638520 1 0 $X=941780 $Y=633100
X1403 4207 2 4200 1 INV1S $T=947360 688920 0 180 $X=946120 $Y=683500
X1404 4171 2 4193 1 INV1S $T=947980 688920 1 180 $X=946740 $Y=688540
X1405 4164 2 4219 1 INV1S $T=950460 557880 1 0 $X=950460 $Y=552460
X1406 4218 2 4210 1 INV1S $T=951700 678840 1 180 $X=950460 $Y=678460
X1407 4196 2 4216 1 INV1S $T=951700 688920 1 0 $X=951700 $Y=683500
X1408 4227 2 4222 1 INV1S $T=953560 678840 1 180 $X=952320 $Y=678460
X1409 600 2 4185 1 INV1S $T=955420 658680 1 0 $X=955420 $Y=653260
X1410 4220 2 4229 1 INV1S $T=958520 557880 1 0 $X=958520 $Y=552460
X1411 4251 2 4259 1 INV1S $T=962240 709080 0 0 $X=962240 $Y=708700
X1412 4272 2 4270 1 INV1S $T=965340 557880 0 180 $X=964100 $Y=552460
X1413 612 2 4280 1 INV1S $T=969680 719160 0 180 $X=968440 $Y=713740
X1414 4280 2 4269 1 INV1S $T=970920 709080 0 180 $X=969680 $Y=703660
X1415 4298 2 4285 1 INV1S $T=972160 678840 1 180 $X=970920 $Y=678460
X1416 615 2 4305 1 INV1S $T=976500 547800 0 180 $X=975260 $Y=542380
X1417 617 2 4303 1 INV1S $T=977120 719160 1 0 $X=977120 $Y=713740
X1418 4303 2 4315 1 INV1S $T=979600 719160 0 180 $X=978360 $Y=713740
X1419 4317 2 4319 1 INV1S $T=978980 618360 1 0 $X=978980 $Y=612940
X1420 4326 2 4327 1 INV1S $T=983940 678840 0 180 $X=982700 $Y=673420
X1421 626 2 4352 1 INV1S $T=990760 699000 1 0 $X=990760 $Y=693580
X1422 4350 2 4364 1 INV1S $T=993240 699000 1 0 $X=993240 $Y=693580
X1423 4362 2 4351 1 INV1S $T=997580 638520 1 180 $X=996340 $Y=638140
X1424 629 2 4376 1 INV1S $T=998200 709080 0 0 $X=998200 $Y=708700
X1425 4357 2 4375 1 INV1S $T=1000680 628440 0 180 $X=999440 $Y=623020
X1426 634 2 4382 1 INV1S $T=1001920 719160 0 180 $X=1000680 $Y=713740
X1427 4396 2 4370 1 INV1S $T=1002540 618360 0 180 $X=1001300 $Y=612940
X1428 4401 2 4393 1 INV1S $T=1004400 719160 0 180 $X=1003160 $Y=713740
X1429 4397 2 4371 1 INV1S $T=1005020 709080 0 180 $X=1003780 $Y=703660
X1430 4408 2 4392 1 INV1S $T=1006880 618360 1 180 $X=1005640 $Y=617980
X1431 4416 2 4381 1 INV1S $T=1008120 699000 0 180 $X=1006880 $Y=693580
X1432 4417 2 640 1 INV1S $T=1014320 547800 0 180 $X=1013080 $Y=542380
X1433 645 2 4395 1 INV1S $T=1018040 699000 1 180 $X=1016800 $Y=698620
X1434 4439 2 4374 1 INV1S $T=1024860 598200 1 180 $X=1023620 $Y=597820
X1435 4454 2 4473 1 INV1S $T=1034160 557880 1 0 $X=1034160 $Y=552460
X1436 4489 2 4483 1 INV1S $T=1045320 557880 0 180 $X=1044080 $Y=552460
X1437 4515 2 4503 1 INV1S $T=1058960 618360 1 180 $X=1057720 $Y=617980
X1438 4537 2 4532 1 INV1S $T=1068880 567960 0 0 $X=1068880 $Y=567580
X1439 701 703 711 718 2 1 MXL2HS $T=265360 567960 0 0 $X=265360 $Y=567580
X1440 769 764 744 757 2 1 MXL2HS $T=286440 567960 1 180 $X=280860 $Y=567580
X1441 713 758 761 725 2 1 MXL2HS $T=280860 608280 0 0 $X=280860 $Y=607900
X1442 836 843 821 830 2 1 MXL2HS $T=300700 578040 1 0 $X=300700 $Y=572620
X1443 930 901 831 894 2 1 MXL2HS $T=316820 608280 1 180 $X=311240 $Y=607900
X1444 993 981 996 961 2 1 MXL2HS $T=327360 608280 0 0 $X=327360 $Y=607900
X1445 1013 1015 1028 1042 2 1 MXL2HS $T=331080 598200 1 0 $X=331080 $Y=592780
X1446 1298 1173 1146 1276 2 1 MXL2HS $T=380680 628440 0 180 $X=375100 $Y=623020
X1447 1414 1412 1402 1396 2 1 MXL2HS $T=403620 567960 1 180 $X=398040 $Y=567580
X1448 93 1419 1451 1431 2 1 MXL2HS $T=413540 557880 0 180 $X=407960 $Y=552460
X1449 1446 1412 1456 1458 2 1 MXL2HS $T=407960 567960 1 0 $X=407960 $Y=562540
X1450 1396 1412 1485 1490 2 1 MXL2HS $T=412920 578040 0 0 $X=412920 $Y=577660
X1451 97 1419 1498 1495 2 1 MXL2HS $T=415400 557880 1 0 $X=415400 $Y=552460
X1452 1431 1412 1470 1511 2 1 MXL2HS $T=417260 567960 0 0 $X=417260 $Y=567580
X1453 1458 1412 1512 1520 2 1 MXL2HS $T=419120 578040 0 0 $X=419120 $Y=577660
X1454 1495 1525 1537 1553 2 1 MXL2HS $T=427180 567960 0 0 $X=427180 $Y=567580
X1455 120 1590 1528 1576 2 1 MXL2HS $T=440200 557880 0 180 $X=434620 $Y=552460
X1456 1576 1525 1594 1603 2 1 MXL2HS $T=435860 567960 0 0 $X=435860 $Y=567580
X1457 1588 124 1524 119 2 1 MXL2HS $T=443920 547800 1 180 $X=438340 $Y=547420
X1458 119 124 1609 1517 2 1 MXL2HS $T=447640 547800 0 180 $X=442060 $Y=542380
X1459 127 1590 1621 1618 2 1 MXL2HS $T=447640 557880 0 180 $X=442060 $Y=552460
X1460 1618 1525 1624 1638 2 1 MXL2HS $T=443300 578040 1 0 $X=443300 $Y=572620
X1461 1660 1590 1643 1588 2 1 MXL2HS $T=453840 547800 1 180 $X=448260 $Y=547420
X1462 129 1590 1644 1661 2 1 MXL2HS $T=448260 557880 1 0 $X=448260 $Y=552460
X1463 1661 1525 1645 1688 2 1 MXL2HS $T=454460 567960 1 0 $X=454460 $Y=562540
X1464 153 149 1755 1778 2 1 MXL2HS $T=480500 709080 1 180 $X=474920 $Y=708700
X1465 150 1684 1794 148 2 1 MXL2HS $T=482360 547800 0 180 $X=476780 $Y=542380
X1466 1823 1684 1800 150 2 1 MXL2HS $T=483600 547800 1 180 $X=478020 $Y=547420
X1467 1787 1797 1801 1770 2 1 MXL2HS $T=483600 648600 0 180 $X=478020 $Y=643180
X1468 1770 1797 1811 1788 2 1 MXL2HS $T=478020 658680 1 0 $X=478020 $Y=653260
X1469 1835 1684 1813 1660 2 1 MXL2HS $T=486080 557880 1 180 $X=480500 $Y=557500
X1470 155 1822 1804 1843 2 1 MXL2HS $T=481120 668760 0 0 $X=481120 $Y=668380
X1471 154 1822 1802 1847 2 1 MXL2HS $T=481740 668760 1 0 $X=481740 $Y=663340
X1472 157 1839 1761 1856 2 1 MXL2HS $T=484220 709080 1 0 $X=484220 $Y=703660
X1473 1778 1822 1805 1864 2 1 MXL2HS $T=487320 678840 1 0 $X=487320 $Y=673420
X1474 1847 1861 1832 1853 2 1 MXL2HS $T=493520 588120 1 180 $X=487940 $Y=587740
X1475 159 1822 1803 1868 2 1 MXL2HS $T=487940 678840 0 0 $X=487940 $Y=678460
X1476 1856 1797 1866 1875 2 1 MXL2HS $T=489180 648600 0 0 $X=489180 $Y=648220
X1477 156 1839 1846 1876 2 1 MXL2HS $T=489180 699000 1 0 $X=489180 $Y=693580
X1478 1853 1861 1837 1823 2 1 MXL2HS $T=495380 588120 0 180 $X=489800 $Y=582700
X1479 162 1797 1872 1860 2 1 MXL2HS $T=489800 648600 1 0 $X=489800 $Y=643180
X1480 164 1839 1834 1879 2 1 MXL2HS $T=490420 709080 0 0 $X=490420 $Y=708700
X1481 158 1839 1867 1901 2 1 MXL2HS $T=494760 699000 0 0 $X=494760 $Y=698620
X1482 1903 1861 1862 1835 2 1 MXL2HS $T=500960 588120 1 180 $X=495380 $Y=587740
X1483 1875 1902 1871 172 2 1 MXL2HS $T=501580 567960 1 180 $X=496000 $Y=567580
X1484 1879 1797 1897 1877 2 1 MXL2HS $T=496000 648600 0 0 $X=496000 $Y=648220
X1485 173 149 1899 1889 2 1 MXL2HS $T=496000 709080 0 0 $X=496000 $Y=708700
X1486 1868 1891 1821 1903 2 1 MXL2HS $T=496620 618360 0 0 $X=496620 $Y=617980
X1487 1843 1891 1827 1906 2 1 MXL2HS $T=496620 628440 1 0 $X=496620 $Y=623020
X1488 1860 1893 1833 177 2 1 MXL2HS $T=497240 608280 1 0 $X=497240 $Y=602860
X1489 1864 1891 1904 1910 2 1 MXL2HS $T=497860 608280 0 0 $X=497860 $Y=607900
X1490 1915 1684 1888 174 2 1 MXL2HS $T=504680 557880 0 180 $X=499100 $Y=552460
X1491 178 1880 1905 1898 2 1 MXL2HS $T=504680 688920 1 180 $X=499100 $Y=688540
X1492 1877 1902 1844 179 2 1 MXL2HS $T=499720 567960 1 0 $X=499720 $Y=562540
X1493 1889 1880 1912 1918 2 1 MXL2HS $T=499720 678840 0 0 $X=499720 $Y=678460
X1494 1908 1902 1909 1915 2 1 MXL2HS $T=500960 588120 1 0 $X=500960 $Y=582700
X1495 1898 1854 1919 1908 2 1 MXL2HS $T=502200 648600 0 0 $X=502200 $Y=648220
X1496 1901 1893 1929 1922 2 1 MXL2HS $T=503440 628440 1 0 $X=503440 $Y=623020
X1497 176 1854 1925 1928 2 1 MXL2HS $T=503440 668760 0 0 $X=503440 $Y=668380
X1498 1926 1902 1921 187 2 1 MXL2HS $T=505920 557880 0 0 $X=505920 $Y=557500
X1499 1876 1893 1917 1939 2 1 MXL2HS $T=505920 618360 1 0 $X=505920 $Y=612940
X1500 1928 1934 1923 1949 2 1 MXL2HS $T=507160 598200 0 0 $X=507160 $Y=597820
X1501 1950 1946 1936 1935 2 1 MXL2HS $T=513360 678840 0 180 $X=507780 $Y=673420
X1502 192 190 185 1937 2 1 MXL2HS $T=513980 719160 0 180 $X=508400 $Y=713740
X1503 1943 191 1933 186 2 1 MXL2HS $T=515220 557880 0 180 $X=509640 $Y=552460
X1504 1961 1938 1951 1943 2 1 MXL2HS $T=515840 567960 0 180 $X=510260 $Y=562540
X1505 1918 1893 1916 1966 2 1 MXL2HS $T=511500 608280 1 0 $X=511500 $Y=602860
X1506 1937 1954 1965 1960 2 1 MXL2HS $T=511500 648600 1 0 $X=511500 $Y=643180
X1507 181 1968 1957 1950 2 1 MXL2HS $T=517700 709080 0 180 $X=512120 $Y=703660
X1508 1906 1934 1953 1958 2 1 MXL2HS $T=518940 598200 1 180 $X=513360 $Y=597820
X1509 1945 1946 1967 1926 2 1 MXL2HS $T=519560 678840 0 180 $X=513980 $Y=673420
X1510 195 1940 1947 1945 2 1 MXL2HS $T=514600 688920 0 0 $X=514600 $Y=688540
X1511 202 1959 1973 1972 2 1 MXL2HS $T=520800 658680 1 180 $X=515220 $Y=658300
X1512 1990 1954 1975 1974 2 1 MXL2HS $T=521420 648600 1 180 $X=515840 $Y=648220
X1513 1935 1996 1964 1978 2 1 MXL2HS $T=522660 618360 0 180 $X=517080 $Y=612940
X1514 200 1968 1969 1979 2 1 MXL2HS $T=517700 709080 1 0 $X=517700 $Y=703660
X1515 1910 1996 1991 1985 2 1 MXL2HS $T=523900 608280 0 180 $X=518320 $Y=602860
X1516 1987 2004 1980 203 2 1 MXL2HS $T=525140 557880 1 180 $X=519560 $Y=557500
X1517 1974 2004 1999 204 2 1 MXL2HS $T=525140 578040 0 180 $X=519560 $Y=572620
X1518 1998 1954 2005 1961 2 1 MXL2HS $T=520180 648600 1 0 $X=520180 $Y=643180
X1519 210 1940 2001 1990 2 1 MXL2HS $T=526380 688920 1 180 $X=520800 $Y=688540
X1520 1960 1959 1981 207 2 1 MXL2HS $T=521420 628440 0 0 $X=521420 $Y=628060
X1521 1972 1996 2015 213 2 1 MXL2HS $T=523280 618360 1 0 $X=523280 $Y=612940
X1522 1997 1934 2027 1992 2 1 MXL2HS $T=525760 608280 0 0 $X=525760 $Y=607900
X1523 1979 1946 2030 2013 2 1 MXL2HS $T=525760 668760 0 0 $X=525760 $Y=668380
X1524 2010 1959 2024 1997 2 1 MXL2HS $T=531960 658680 1 180 $X=526380 $Y=658300
X1525 1982 2028 2023 1987 2 1 MXL2HS $T=527000 638520 1 0 $X=527000 $Y=633100
X1526 2000 1959 2037 1982 2 1 MXL2HS $T=527620 648600 1 0 $X=527620 $Y=643180
X1527 219 1940 2011 1998 2 1 MXL2HS $T=533200 688920 1 180 $X=527620 $Y=688540
X1528 2013 1996 2040 222 2 1 MXL2HS $T=529480 618360 1 0 $X=529480 $Y=612940
X1529 1966 1938 2020 2019 2 1 MXL2HS $T=530100 578040 0 0 $X=530100 $Y=577660
X1530 201 2039 2045 2048 2 1 MXL2HS $T=530100 699000 0 0 $X=530100 $Y=698620
X1531 227 226 220 2000 2 1 MXL2HS $T=537540 719160 0 180 $X=531960 $Y=713740
X1532 223 1940 2061 2063 2 1 MXL2HS $T=533200 688920 0 0 $X=533200 $Y=688540
X1533 1922 1996 2054 2032 2 1 MXL2HS $T=539400 608280 1 180 $X=533820 $Y=607900
X1534 224 1946 2038 2068 2 1 MXL2HS $T=534440 678840 1 0 $X=534440 $Y=673420
X1535 1978 191 2066 2073 2 1 MXL2HS $T=535060 547800 0 0 $X=535060 $Y=547420
X1536 1949 1938 2070 2003 2 1 MXL2HS $T=536300 578040 0 0 $X=536300 $Y=577660
X1537 217 2039 2065 2010 2 1 MXL2HS $T=536300 709080 1 0 $X=536300 $Y=703660
X1538 1992 1938 2078 231 2 1 MXL2HS $T=536920 557880 0 0 $X=536920 $Y=557500
X1539 2063 2041 2079 233 2 1 MXL2HS $T=537540 658680 0 0 $X=537540 $Y=658300
X1540 2087 226 2075 208 2 1 MXL2HS $T=543740 719160 0 180 $X=538160 $Y=713740
X1541 228 2039 2089 2093 2 1 MXL2HS $T=539400 699000 0 0 $X=539400 $Y=698620
X1542 2033 2081 2071 2095 2 1 MXL2HS $T=540020 608280 0 0 $X=540020 $Y=607900
X1543 2048 2041 2092 2084 2 1 MXL2HS $T=541260 658680 1 0 $X=541260 $Y=653260
X1544 2068 2028 2098 2094 2 1 MXL2HS $T=543120 628440 0 0 $X=543120 $Y=628060
X1545 2093 2041 2097 2033 2 1 MXL2HS $T=549320 678840 0 180 $X=543740 $Y=673420
X1546 235 2039 2101 2103 2 1 MXL2HS $T=544360 709080 1 0 $X=544360 $Y=703660
X1547 1939 2081 2109 2036 2 1 MXL2HS $T=546220 608280 0 0 $X=546220 $Y=607900
X1548 2103 2041 2113 2050 2 1 MXL2HS $T=546840 668760 0 0 $X=546840 $Y=668380
X1549 2111 2028 2106 2043 2 1 MXL2HS $T=549320 628440 0 0 $X=549320 $Y=628060
X1550 2130 2125 2100 2080 2 1 MXL2HS $T=557380 648600 1 180 $X=551800 $Y=648220
X1551 2095 2081 2119 2131 2 1 MXL2HS $T=552420 608280 0 0 $X=552420 $Y=607900
X1552 251 2090 2120 2111 2 1 MXL2HS $T=558000 688920 1 180 $X=552420 $Y=688540
X1553 2036 2051 2136 2141 2 1 MXL2HS $T=554280 608280 1 0 $X=554280 $Y=602860
X1554 240 2090 2137 2130 2 1 MXL2HS $T=554280 678840 0 0 $X=554280 $Y=678460
X1555 2050 2051 2142 2128 2 1 MXL2HS $T=556140 588120 0 0 $X=556140 $Y=587740
X1556 2153 2125 2121 2132 2 1 MXL2HS $T=561720 668760 0 180 $X=556140 $Y=663340
X1557 2154 2039 2138 2087 2 1 MXL2HS $T=561720 709080 0 180 $X=556140 $Y=703660
X1558 2080 2150 2139 2116 2 1 MXL2HS $T=562960 618360 1 180 $X=557380 $Y=617980
X1559 2159 2039 2144 254 2 1 MXL2HS $T=562960 699000 1 180 $X=557380 $Y=698620
X1560 2084 2147 2155 2124 2 1 MXL2HS $T=558620 557880 1 0 $X=558620 $Y=552460
X1561 2043 2147 2135 2133 2 1 MXL2HS $T=559240 567960 1 0 $X=559240 $Y=562540
X1562 2149 2125 2156 2165 2 1 MXL2HS $T=559240 648600 0 0 $X=559240 $Y=648220
X1563 2132 2125 2134 2149 2 1 MXL2HS $T=559240 658680 1 0 $X=559240 $Y=653260
X1564 2019 2051 2168 2173 2 1 MXL2HS $T=561720 588120 0 0 $X=561720 $Y=587740
X1565 2094 2147 2170 257 2 1 MXL2HS $T=562340 557880 0 0 $X=562340 $Y=557500
X1566 1958 2051 2129 2177 2 1 MXL2HS $T=562340 598200 0 0 $X=562340 $Y=597820
X1567 258 2090 2152 2153 2 1 MXL2HS $T=567920 678840 1 180 $X=562340 $Y=678460
X1568 2116 2150 2161 2188 2 1 MXL2HS $T=564820 618360 0 0 $X=564820 $Y=617980
X1569 257 2147 2180 2191 2 1 MXL2HS $T=565440 557880 1 0 $X=565440 $Y=552460
X1570 2194 2125 2181 2175 2 1 MXL2HS $T=571020 658680 0 180 $X=565440 $Y=653260
X1571 2032 2174 2171 2197 2 1 MXL2HS $T=566680 608280 1 0 $X=566680 $Y=602860
X1572 2175 2125 2189 2176 2 1 MXL2HS $T=573500 668760 0 180 $X=567920 $Y=663340
X1573 2176 2090 2190 2159 2 1 MXL2HS $T=573500 678840 1 180 $X=567920 $Y=678460
X1574 2212 2090 2199 2154 2 1 MXL2HS $T=577220 688920 1 180 $X=571640 $Y=688540
X1575 2124 2147 2213 2218 2 1 MXL2HS $T=573500 557880 0 0 $X=573500 $Y=557500
X1576 1985 2174 2216 2219 2 1 MXL2HS $T=573500 608280 1 0 $X=573500 $Y=602860
X1577 2227 2090 2183 2212 2 1 MXL2HS $T=580320 678840 0 180 $X=574740 $Y=673420
X1578 2003 2214 2222 2229 2 1 MXL2HS $T=575360 588120 1 0 $X=575360 $Y=582700
X1579 262 264 2160 267 2 1 MXL2HS $T=575980 547800 1 0 $X=575980 $Y=542380
X1580 203 2214 2166 2236 2 1 MXL2HS $T=577840 567960 0 0 $X=577840 $Y=567580
X1581 2238 2235 2205 263 2 1 MXL2HS $T=584040 709080 1 180 $X=578460 $Y=708700
X1582 2241 2235 2208 268 2 1 MXL2HS $T=585280 699000 1 180 $X=579700 $Y=698620
X1583 2219 2150 2215 2247 2 1 MXL2HS $T=580940 618360 1 0 $X=580940 $Y=612940
X1584 270 264 2224 2248 2 1 MXL2HS $T=581560 547800 1 0 $X=581560 $Y=542380
X1585 2128 2214 2244 2249 2 1 MXL2HS $T=581560 588120 1 0 $X=581560 $Y=582700
X1586 2177 2150 2231 2253 2 1 MXL2HS $T=582800 628440 1 0 $X=582800 $Y=623020
X1587 2256 2252 2228 2227 2 1 MXL2HS $T=589000 658680 0 180 $X=583420 $Y=653260
X1588 2250 272 2232 2238 2 1 MXL2HS $T=589000 688920 1 180 $X=583420 $Y=688540
X1589 2133 2214 2225 2260 2 1 MXL2HS $T=584040 567960 0 0 $X=584040 $Y=567580
X1590 2268 2252 2240 2250 2 1 MXL2HS $T=590860 668760 0 180 $X=585280 $Y=663340
X1591 234 2258 2243 2277 2 1 MXL2HS $T=587140 557880 1 0 $X=587140 $Y=552460
X1592 2280 2235 2263 274 2 1 MXL2HS $T=592720 709080 0 180 $X=587140 $Y=703660
X1593 2281 2235 2245 2241 2 1 MXL2HS $T=593960 699000 1 180 $X=588380 $Y=698620
X1594 2267 2252 2265 2288 2 1 MXL2HS $T=589000 658680 1 0 $X=589000 $Y=653260
X1595 2131 2282 2294 2295 2 1 MXL2HS $T=590860 618360 1 0 $X=590860 $Y=612940
X1596 2247 2252 2269 2299 2 1 MXL2HS $T=591480 648600 1 0 $X=591480 $Y=643180
X1597 2253 2282 2291 2267 2 1 MXL2HS $T=592100 628440 1 0 $X=592100 $Y=623020
X1598 2300 2252 2292 2281 2 1 MXL2HS $T=597680 668760 1 180 $X=592100 $Y=668380
X1599 2073 2258 2275 2303 2 1 MXL2HS $T=592720 547800 0 0 $X=592720 $Y=547420
X1600 2296 2252 2305 2309 2 1 MXL2HS $T=594580 648600 0 0 $X=594580 $Y=648220
X1601 2311 2235 2302 2280 2 1 MXL2HS $T=600780 699000 1 180 $X=595200 $Y=698620
X1602 284 2319 2310 278 2 1 MXL2HS $T=603260 719160 0 180 $X=597680 $Y=713740
X1603 279 2258 2274 285 2 1 MXL2HS $T=598300 547800 0 0 $X=598300 $Y=547420
X1604 2197 2282 2287 2296 2 1 MXL2HS $T=603880 618360 0 180 $X=598300 $Y=612940
X1605 231 2312 2314 2331 2 1 MXL2HS $T=598920 567960 1 0 $X=598920 $Y=562540
X1606 2295 2306 2329 2334 2 1 MXL2HS $T=599540 648600 1 0 $X=599540 $Y=643180
X1607 2188 2282 2234 2328 2 1 MXL2HS $T=601400 628440 1 0 $X=601400 $Y=623020
X1608 2288 2330 2308 2342 2 1 MXL2HS $T=602020 678840 0 0 $X=602020 $Y=678460
X1609 2249 2337 2289 2349 2 1 MXL2HS $T=603880 588120 1 0 $X=603880 $Y=582700
X1610 2173 2337 2284 2350 2 1 MXL2HS $T=603880 598200 1 0 $X=603880 $Y=592780
X1611 2354 2330 2301 284 2 1 MXL2HS $T=610080 699000 0 180 $X=604500 $Y=693580
X1612 288 2312 2343 2355 2 1 MXL2HS $T=605120 547800 0 0 $X=605120 $Y=547420
X1613 2218 2312 2335 2356 2 1 MXL2HS $T=605120 567960 1 0 $X=605120 $Y=562540
X1614 2340 2306 2347 2357 2 1 MXL2HS $T=605120 648600 1 0 $X=605120 $Y=643180
X1615 2141 2282 2339 2340 2 1 MXL2HS $T=611320 618360 0 180 $X=605740 $Y=612940
X1616 2342 2319 2333 289 2 1 MXL2HS $T=611940 709080 0 180 $X=606360 $Y=703660
X1617 2309 2364 2348 2354 2 1 MXL2HS $T=614420 678840 1 180 $X=608840 $Y=678460
X1618 2373 2330 2359 2311 2 1 MXL2HS $T=615040 688920 1 180 $X=609460 $Y=688540
X1619 2328 2306 2374 2378 2 1 MXL2HS $T=610700 638520 1 0 $X=610700 $Y=633100
X1620 2299 2364 2380 2384 2 1 MXL2HS $T=611940 668760 1 0 $X=611940 $Y=663340
X1621 2236 2386 2313 2372 2 1 MXL2HS $T=618760 578040 0 180 $X=613180 $Y=572620
X1622 2277 2312 2385 2396 2 1 MXL2HS $T=614420 567960 1 0 $X=614420 $Y=562540
X1623 2334 2364 2367 2399 2 1 MXL2HS $T=615040 658680 0 0 $X=615040 $Y=658300
X1624 2399 2319 2365 294 2 1 MXL2HS $T=621240 699000 1 180 $X=615660 $Y=698620
X1625 2350 2387 2397 2403 2 1 MXL2HS $T=616280 618360 0 0 $X=616280 $Y=617980
X1626 267 2376 286 2408 2 1 MXL2HS $T=616900 547800 1 0 $X=616900 $Y=542380
X1627 2229 2337 2370 2390 2 1 MXL2HS $T=622480 588120 1 180 $X=616900 $Y=587740
X1628 2357 2364 2401 2409 2 1 MXL2HS $T=616900 678840 0 0 $X=616900 $Y=678460
X1629 2349 2387 2398 2412 2 1 MXL2HS $T=617520 628440 1 0 $X=617520 $Y=623020
X1630 2415 2319 2388 299 2 1 MXL2HS $T=625580 719160 0 180 $X=620000 $Y=713740
X1631 2260 2386 2393 2411 2 1 MXL2HS $T=620620 578040 0 0 $X=620620 $Y=577660
X1632 2411 2337 2395 2427 2 1 MXL2HS $T=621240 608280 1 0 $X=621240 $Y=602860
X1633 2378 2364 2426 2415 2 1 MXL2HS $T=622480 678840 0 0 $X=622480 $Y=678460
X1634 285 2376 301 2432 2 1 MXL2HS $T=623100 547800 1 0 $X=623100 $Y=542380
X1635 2438 2422 2450 2373 2 1 MXL2HS $T=627440 638520 1 0 $X=627440 $Y=633100
X1636 2412 2422 2383 2443 2 1 MXL2HS $T=627440 638520 0 0 $X=627440 $Y=638140
X1637 2443 2444 2453 307 2 1 MXL2HS $T=628060 699000 0 0 $X=628060 $Y=698620
X1638 2331 2386 2454 2430 2 1 MXL2HS $T=628680 588120 1 0 $X=628680 $Y=582700
X1639 2409 303 2457 308 2 1 MXL2HS $T=628680 719160 1 0 $X=628680 $Y=713740
X1640 2390 2387 2467 2438 2 1 MXL2HS $T=631780 618360 0 0 $X=631780 $Y=617980
X1641 2191 2405 2445 2473 2 1 MXL2HS $T=632400 567960 1 0 $X=632400 $Y=562540
X1642 2403 2422 2419 2464 2 1 MXL2HS $T=638600 638520 1 180 $X=633020 $Y=638140
X1643 2372 2337 2407 2474 2 1 MXL2HS $T=633640 598200 0 0 $X=633640 $Y=597820
X1644 2427 2404 2414 2477 2 1 MXL2HS $T=633640 668760 1 0 $X=633640 $Y=663340
X1645 2303 2386 2446 2478 2 1 MXL2HS $T=634260 567960 0 0 $X=634260 $Y=567580
X1646 2477 2444 2456 310 2 1 MXL2HS $T=639840 699000 1 180 $X=634260 $Y=698620
X1647 2430 2337 2460 2476 2 1 MXL2HS $T=634880 598200 1 0 $X=634880 $Y=592780
X1648 2248 2471 2479 2485 2 1 MXL2HS $T=636120 557880 1 0 $X=636120 $Y=552460
X1649 1520 2386 2481 315 2 1 MXL2HS $T=636740 578040 0 0 $X=636740 $Y=577660
X1650 2384 303 2475 313 2 1 MXL2HS $T=642320 709080 1 180 $X=636740 $Y=708700
X1651 2464 2488 2452 314 2 1 MXL2HS $T=642940 688920 0 180 $X=637360 $Y=683500
X1652 309 2471 316 2501 2 1 MXL2HS $T=639220 547800 0 0 $X=639220 $Y=547420
X1653 2432 2472 2482 2502 2 1 MXL2HS $T=639220 608280 1 0 $X=639220 $Y=602860
X1654 2474 2484 2493 2268 2 1 MXL2HS $T=639220 648600 0 0 $X=639220 $Y=648220
X1655 2476 2404 2496 2487 2 1 MXL2HS $T=639840 668760 1 0 $X=639840 $Y=663340
X1656 2487 2444 2500 319 2 1 MXL2HS $T=639840 699000 0 0 $X=639840 $Y=698620
X1657 1553 2405 2491 320 2 1 MXL2HS $T=641700 567960 0 0 $X=641700 $Y=567580
X1658 2408 2509 2480 2498 2 1 MXL2HS $T=647280 618360 1 180 $X=641700 $Y=617980
X1659 2355 2472 2470 2503 2 1 MXL2HS $T=648520 618360 0 180 $X=642940 $Y=612940
X1660 2503 2484 2507 2300 2 1 MXL2HS $T=648520 658680 0 180 $X=642940 $Y=653260
X1661 2511 2488 2497 318 2 1 MXL2HS $T=649140 688920 0 180 $X=643560 $Y=683500
X1662 2502 2404 2495 2511 2 1 MXL2HS $T=651000 668760 0 180 $X=645420 $Y=663340
X1663 2522 2520 2512 322 2 1 MXL2HS $T=651620 699000 0 180 $X=646040 $Y=693580
X1664 2485 2472 2528 2535 2 1 MXL2HS $T=647900 608280 1 0 $X=647900 $Y=602860
X1665 1788 2405 2527 2539 2 1 MXL2HS $T=648520 567960 0 0 $X=648520 $Y=567580
X1666 2542 327 2524 2516 2 1 MXL2HS $T=654720 547800 1 180 $X=649140 $Y=547420
X1667 2535 2484 2489 2194 2 1 MXL2HS $T=654720 648600 0 180 $X=649140 $Y=643180
X1668 1688 2526 2541 328 2 1 MXL2HS $T=650380 567960 1 0 $X=650380 $Y=562540
X1669 1490 2526 2544 2534 2 1 MXL2HS $T=650380 578040 0 0 $X=650380 $Y=577660
X1670 2473 2509 2514 2550 2 1 MXL2HS $T=650380 628440 0 0 $X=650380 $Y=628060
X1671 2534 327 2547 2542 2 1 MXL2HS $T=651620 557880 1 0 $X=651620 $Y=552460
X1672 2396 2509 2548 2556 2 1 MXL2HS $T=651620 618360 1 0 $X=651620 $Y=612940
X1673 2540 2404 2552 2543 2 1 MXL2HS $T=652240 668760 1 0 $X=652240 $Y=663340
X1674 2356 2509 2537 2540 2 1 MXL2HS $T=652860 628440 1 0 $X=652860 $Y=623020
X1675 2543 2488 2555 330 2 1 MXL2HS $T=652860 688920 1 0 $X=652860 $Y=683500
X1676 2501 2472 2559 2568 2 1 MXL2HS $T=654720 608280 1 0 $X=654720 $Y=602860
X1677 2556 2484 2560 2256 2 1 MXL2HS $T=661540 648600 0 180 $X=655960 $Y=643180
X1678 1638 2526 2558 334 2 1 MXL2HS $T=656580 578040 1 0 $X=656580 $Y=572620
X1679 2498 2484 2572 2530 2 1 MXL2HS $T=656580 638520 0 0 $X=656580 $Y=638140
X1680 2550 2484 2564 2522 2 1 MXL2HS $T=662160 648600 1 180 $X=656580 $Y=648220
X1681 2583 327 2567 2575 2 1 MXL2HS $T=665260 557880 1 180 $X=659680 $Y=557500
X1682 2478 2509 2574 2577 2 1 MXL2HS $T=659680 628440 1 0 $X=659680 $Y=623020
X1683 2551 2520 2561 333 2 1 MXL2HS $T=665260 699000 1 180 $X=659680 $Y=698620
X1684 2577 2580 2587 2570 2 1 MXL2HS $T=662160 658680 0 0 $X=662160 $Y=658300
X1685 2530 2520 2592 2595 2 1 MXL2HS $T=665260 699000 0 0 $X=665260 $Y=698620
X1686 2539 327 2601 2583 2 1 MXL2HS $T=668360 557880 0 0 $X=668360 $Y=557500
X1687 2570 2520 2585 338 2 1 MXL2HS $T=674560 699000 0 180 $X=668980 $Y=693580
X1688 2597 340 2578 2605 2 1 MXL2HS $T=669600 547800 0 0 $X=669600 $Y=547420
X1689 2568 2580 2591 2551 2 1 MXL2HS $T=675180 668760 0 180 $X=669600 $Y=663340
X1690 1603 2526 2607 346 2 1 MXL2HS $T=671460 567960 1 0 $X=671460 $Y=562540
X1691 1511 2526 2590 2597 2 1 MXL2HS $T=671460 578040 0 0 $X=671460 $Y=577660
X1692 2516 342 2610 347 2 1 MXL2HS $T=671460 719160 1 0 $X=671460 $Y=713740
X1693 345 2580 2619 350 2 1 MXL2HS $T=674560 699000 1 0 $X=674560 $Y=693580
X1694 2595 342 2586 351 2 1 MXL2HS $T=676420 709080 0 0 $X=676420 $Y=708700
X1695 348 2580 2623 352 2 1 MXL2HS $T=677040 699000 0 0 $X=677040 $Y=698620
X1696 2605 340 2625 2617 2 1 MXL2HS $T=678280 547800 0 0 $X=678280 $Y=547420
X1697 2617 2580 2632 354 2 1 MXL2HS $T=678900 678840 1 0 $X=678900 $Y=673420
X1698 2575 2580 2616 355 2 1 MXL2HS $T=679520 688920 1 0 $X=679520 $Y=683500
X1699 2924 2916 2936 2950 2 1 MXL2HS $T=727260 557880 0 0 $X=727260 $Y=557500
X1700 3377 3380 442 3382 2 1 MXL2HS $T=795460 567960 0 0 $X=795460 $Y=567580
X1701 3528 3498 467 3522 2 1 MXL2HS $T=821500 598200 0 0 $X=821500 $Y=597820
X1702 4298 4289 4267 4285 2 1 MXL2HS $T=974020 678840 0 180 $X=968440 $Y=673420
X1703 4315 4311 4306 4303 2 1 MXL2HS $T=979600 678840 1 180 $X=974020 $Y=678460
X1704 4350 4347 4361 4364 2 1 MXL2HS $T=990140 688920 0 0 $X=990140 $Y=688540
X1705 4376 633 4368 4371 2 1 MXL2HS $T=1001920 709080 0 180 $X=996340 $Y=703660
X1706 4375 631 4346 4392 2 1 MXL2HS $T=998820 618360 0 0 $X=998820 $Y=617980
X1707 4381 633 4355 4395 2 1 MXL2HS $T=1000060 699000 1 0 $X=1000060 $Y=693580
X1708 4382 633 4391 4393 2 1 MXL2HS $T=1000060 709080 0 0 $X=1000060 $Y=708700
X1709 4473 631 4445 4483 2 1 MXL2HS $T=1038500 557880 1 0 $X=1038500 $Y=552460
X1710 4491 631 4462 4503 2 1 MXL2HS $T=1045940 618360 0 0 $X=1045940 $Y=617980
X1711 166 161 1 2 INV8 $T=487940 557880 1 0 $X=487940 $Y=552460
X1712 1555 3 1 2 INV12CK $T=432140 598200 0 180 $X=422220 $Y=592780
X1713 1555 11 1 2 INV12CK $T=442060 638520 0 0 $X=442060 $Y=638140
X1714 230 116 1 2 INV12CK $T=540640 547800 0 0 $X=540640 $Y=547420
X1715 269 1791 1 2 INV12CK $T=582180 658680 0 180 $X=572260 $Y=653260
X1716 269 152 1 2 INV12CK $T=580940 668760 0 0 $X=580940 $Y=668380
X1717 230 250 1 2 INV12CK $T=602640 557880 0 180 $X=592720 $Y=552460
X1718 283 2286 1 2 INV12CK $T=602640 709080 0 180 $X=592720 $Y=703660
X1719 269 271 1 2 INV12CK $T=604500 658680 0 180 $X=594580 $Y=653260
X1720 2351 230 1 2 INV12CK $T=611320 608280 0 180 $X=601400 $Y=602860
X1721 2351 269 1 2 INV12CK $T=608220 658680 1 0 $X=608220 $Y=653260
X1722 331 2351 1 2 INV12CK $T=657820 668760 0 0 $X=657820 $Y=668380
X1723 2286 331 1 2 INV12CK $T=657820 678840 0 0 $X=657820 $Y=678460
X1724 2614 2290 1 2 INV12CK $T=703080 658680 0 180 $X=693160 $Y=653260
X1725 2614 465 1 2 INV12CK $T=829560 658680 0 180 $X=819640 $Y=653260
X1726 2286 523 1 2 INV12CK $T=880400 547800 0 0 $X=880400 $Y=547420
X1727 4399 585 1 2 INV12CK $T=1006260 557880 0 0 $X=1006260 $Y=557500
X1728 4394 4080 1 2 INV12CK $T=1013700 598200 0 0 $X=1013700 $Y=597820
X1729 4394 4451 1 2 INV12CK $T=1035400 598200 0 0 $X=1035400 $Y=597820
X1730 4399 650 1 2 INV12CK $T=1055240 557880 0 180 $X=1045320 $Y=552460
X1731 705 685 1 2 692 AN2 $T=266600 578040 1 180 $X=264120 $Y=577660
X1732 1601 1605 1 2 1656 AN2 $T=448880 638520 1 0 $X=448880 $Y=633100
X1733 2700 2711 1 2 2734 AN2 $T=700600 567960 1 0 $X=700600 $Y=562540
X1734 2683 2765 1 2 2747 AN2 $T=708660 608280 0 180 $X=706180 $Y=602860
X1735 2805 2837 1 2 2847 AN2 $T=717340 618360 1 0 $X=717340 $Y=612940
X1736 2858 2781 1 2 2867 AN2 $T=719200 688920 0 0 $X=719200 $Y=688540
X1737 3175 3186 1 2 3195 AN2 $T=766940 658680 1 0 $X=766940 $Y=653260
X1738 3185 3264 1 2 3289 AN2 $T=779960 648600 1 0 $X=779960 $Y=643180
X1739 3501 3400 1 2 3514 AN2 $T=816540 638520 1 0 $X=816540 $Y=633100
X1740 616 614 1 2 4298 AN2 $T=974020 709080 0 180 $X=971540 $Y=703660
X1741 678 681 677 1 2 ND2 $T=259160 638520 0 180 $X=257300 $Y=633100
X1742 737 705 716 1 2 ND2 $T=276520 598200 1 0 $X=276520 $Y=592780
X1743 797 801 747 1 2 ND2 $T=292020 628440 1 180 $X=290160 $Y=628060
X1744 762 782 771 1 2 ND2 $T=290780 608280 0 0 $X=290780 $Y=607900
X1745 801 746 808 1 2 ND2 $T=295120 628440 0 180 $X=293260 $Y=623020
X1746 814 793 839 1 2 ND2 $T=295740 688920 1 0 $X=295740 $Y=683500
X1747 826 830 805 1 2 ND2 $T=298220 598200 1 0 $X=298220 $Y=592780
X1748 817 808 795 1 2 ND2 $T=298220 628440 0 0 $X=298220 $Y=628060
X1749 814 812 854 1 2 ND2 $T=298840 688920 1 0 $X=298840 $Y=683500
X1750 847 855 860 1 2 ND2 $T=301320 598200 1 0 $X=301320 $Y=592780
X1751 854 790 839 1 2 ND2 $T=302560 688920 1 0 $X=302560 $Y=683500
X1752 14 16 8 1 2 ND2 $T=306900 547800 0 180 $X=305040 $Y=542380
X1753 886 805 899 1 2 ND2 $T=308140 598200 0 0 $X=308140 $Y=597820
X1754 18 903 16 1 2 ND2 $T=311860 547800 0 180 $X=310000 $Y=542380
X1755 905 895 871 1 2 ND2 $T=310620 648600 1 0 $X=310620 $Y=643180
X1756 889 915 865 1 2 ND2 $T=313100 547800 1 180 $X=311240 $Y=547420
X1757 913 912 884 1 2 ND2 $T=313720 557880 0 180 $X=311860 $Y=552460
X1758 926 859 948 1 2 ND2 $T=316820 608280 0 0 $X=316820 $Y=607900
X1759 938 948 944 1 2 ND2 $T=320540 608280 1 0 $X=320540 $Y=602860
X1760 851 970 934 1 2 ND2 $T=323640 638520 0 180 $X=321780 $Y=633100
X1761 940 979 909 1 2 ND2 $T=324880 567960 0 180 $X=323020 $Y=562540
X1762 941 987 967 1 2 ND2 $T=326120 598200 1 0 $X=326120 $Y=592780
X1763 988 999 987 1 2 ND2 $T=327360 588120 0 0 $X=327360 $Y=587740
X1764 990 1003 816 1 2 ND2 $T=329840 547800 0 180 $X=327980 $Y=542380
X1765 1032 1031 973 1 2 ND2 $T=333560 557880 1 180 $X=331700 $Y=557500
X1766 1007 1053 991 1 2 ND2 $T=338520 578040 1 180 $X=336660 $Y=577660
X1767 1048 38 1003 1 2 ND2 $T=337280 547800 1 0 $X=337280 $Y=542380
X1768 1033 1007 1028 1 2 ND2 $T=337900 588120 1 0 $X=337900 $Y=582700
X1769 1058 1030 1047 1 2 ND2 $T=337900 678840 0 0 $X=337900 $Y=678460
X1770 1040 40 1038 1 2 ND2 $T=341000 547800 0 0 $X=341000 $Y=547420
X1771 44 1080 1087 1 2 ND2 $T=344720 719160 1 0 $X=344720 $Y=713740
X1772 943 1114 1041 1 2 ND2 $T=349060 567960 0 180 $X=347200 $Y=562540
X1773 46 1118 1112 1 2 ND2 $T=349680 699000 0 0 $X=349680 $Y=698620
X1774 1060 1100 1112 1 2 ND2 $T=349680 709080 1 0 $X=349680 $Y=703660
X1775 1121 1045 1131 1 2 ND2 $T=350300 628440 0 0 $X=350300 $Y=628060
X1776 1008 1132 1074 1 2 ND2 $T=354020 557880 1 180 $X=352160 $Y=557500
X1777 1160 1161 868 1 2 ND2 $T=357740 648600 0 0 $X=357740 $Y=648220
X1778 1172 1171 1152 1 2 ND2 $T=360220 557880 1 180 $X=358360 $Y=557500
X1779 1147 799 1189 1 2 ND2 $T=360840 638520 0 0 $X=360840 $Y=638140
X1780 1194 1193 1114 1 2 ND2 $T=363940 567960 0 180 $X=362080 $Y=562540
X1781 1113 55 1134 1 2 ND2 $T=364560 547800 0 180 $X=362700 $Y=542380
X1782 1166 1213 1158 1 2 ND2 $T=366420 578040 1 180 $X=364560 $Y=577660
X1783 1170 57 1218 1 2 ND2 $T=365180 547800 1 0 $X=365180 $Y=542380
X1784 1226 1278 1132 1 2 ND2 $T=375100 557880 0 180 $X=373240 $Y=552460
X1785 1185 1283 1264 1 2 ND2 $T=376340 638520 0 180 $X=374480 $Y=633100
X1786 64 1220 1250 1 2 ND2 $T=377580 547800 0 180 $X=375720 $Y=542380
X1787 1262 1310 1316 1 2 ND2 $T=381300 547800 0 0 $X=381300 $Y=547420
X1788 1313 1309 1236 1 2 ND2 $T=381920 618360 0 0 $X=381920 $Y=617980
X1789 1330 1327 1317 1 2 ND2 $T=384400 688920 1 180 $X=382540 $Y=688540
X1790 1327 1275 1318 1 2 ND2 $T=384400 699000 0 180 $X=382540 $Y=693580
X1791 1347 1279 1287 1 2 ND2 $T=387500 588120 0 180 $X=385640 $Y=582700
X1792 1334 1318 1340 1 2 ND2 $T=386880 699000 1 0 $X=386880 $Y=693580
X1793 1374 1325 1360 1 2 ND2 $T=394320 547800 0 0 $X=394320 $Y=547420
X1794 1364 1366 1418 1 2 ND2 $T=401140 678840 0 0 $X=401140 $Y=678460
X1795 1426 1429 1366 1 2 ND2 $T=405480 678840 1 180 $X=403620 $Y=678460
X1796 84 1424 1419 1 2 ND2 $T=406100 547800 1 0 $X=406100 $Y=542380
X1797 1453 1436 1472 1 2 ND2 $T=410440 648600 1 0 $X=410440 $Y=643180
X1798 94 1464 1419 1 2 ND2 $T=413540 547800 1 180 $X=411680 $Y=547420
X1799 1474 1489 1497 1 2 ND2 $T=416640 638520 0 0 $X=416640 $Y=638140
X1800 1494 1488 101 1 2 ND2 $T=417260 709080 0 0 $X=417260 $Y=708700
X1801 1486 1467 1500 1 2 ND2 $T=420980 678840 1 180 $X=419120 $Y=678460
X1802 1534 1544 1493 1 2 ND2 $T=429040 608280 0 180 $X=427180 $Y=602860
X1803 108 1509 1523 1 2 ND2 $T=427180 709080 1 0 $X=427180 $Y=703660
X1804 1613 1629 1632 1 2 ND2 $T=443300 678840 1 0 $X=443300 $Y=673420
X1805 1611 1632 1626 1 2 ND2 $T=445160 688920 0 0 $X=445160 $Y=688540
X1806 1625 1639 1556 1 2 ND2 $T=448260 628440 1 180 $X=446400 $Y=628060
X1807 1450 1705 1669 1 2 ND2 $T=461280 557880 0 180 $X=459420 $Y=552460
X1808 1695 1710 1701 1 2 ND2 $T=463140 578040 0 180 $X=461280 $Y=572620
X1809 1706 1718 1708 1 2 ND2 $T=465000 557880 1 180 $X=463140 $Y=557500
X1810 1729 1715 142 1 2 ND2 $T=466240 618360 0 180 $X=464380 $Y=612940
X1811 1744 1736 1727 1 2 ND2 $T=468720 608280 1 180 $X=466860 $Y=607900
X1812 1735 1748 1712 1 2 ND2 $T=470580 578040 1 180 $X=468720 $Y=577660
X1813 1685 1766 1697 1 2 ND2 $T=470580 588120 0 180 $X=468720 $Y=582700
X1814 1760 1754 1734 1 2 ND2 $T=472440 608280 0 180 $X=470580 $Y=602860
X1815 1772 1756 1730 1 2 ND2 $T=474300 557880 0 180 $X=472440 $Y=552460
X1816 1733 1775 1702 1 2 ND2 $T=474300 598200 0 180 $X=472440 $Y=592780
X1817 1751 1789 1715 1 2 ND2 $T=477400 618360 0 180 $X=475540 $Y=612940
X1818 1769 1814 1736 1 2 ND2 $T=481120 608280 1 180 $X=479260 $Y=607900
X1819 238 1850 2028 1 2 ND2 $T=546840 638520 0 0 $X=546840 $Y=638140
X1820 238 2151 249 1 2 ND2 $T=558000 628440 1 180 $X=556140 $Y=628060
X1821 2626 2638 2615 1 2 ND2 $T=683860 608280 0 180 $X=682000 $Y=602860
X1822 2628 2679 2639 1 2 ND2 $T=690680 618360 0 0 $X=690680 $Y=617980
X1823 2675 2667 2694 1 2 ND2 $T=693160 567960 1 0 $X=693160 $Y=562540
X1824 2682 2690 2679 1 2 ND2 $T=693160 618360 0 0 $X=693160 $Y=617980
X1825 2634 2695 2687 1 2 ND2 $T=695640 608280 1 0 $X=695640 $Y=602860
X1826 2744 2757 2742 1 2 ND2 $T=704320 557880 0 0 $X=704320 $Y=557500
X1827 2757 2768 2756 1 2 ND2 $T=709280 557880 1 180 $X=707420 $Y=557500
X1828 2751 2756 2747 1 2 ND2 $T=707420 567960 1 0 $X=707420 $Y=562540
X1829 2753 2779 2721 1 2 ND2 $T=709280 678840 0 180 $X=707420 $Y=673420
X1830 2771 2752 2746 1 2 ND2 $T=709280 547800 0 0 $X=709280 $Y=547420
X1831 2770 2801 2781 1 2 ND2 $T=711140 699000 1 0 $X=711140 $Y=693580
X1832 2811 2804 2794 1 2 ND2 $T=714240 598200 1 180 $X=712380 $Y=597820
X1833 2818 378 2768 1 2 ND2 $T=714860 547800 1 180 $X=713000 $Y=547420
X1834 2766 2806 2645 1 2 ND2 $T=716100 638520 1 180 $X=714240 $Y=638140
X1835 2766 2832 2792 1 2 ND2 $T=716100 638520 0 0 $X=716100 $Y=638140
X1836 2728 2855 2827 1 2 ND2 $T=718580 588120 1 180 $X=716720 $Y=587740
X1837 2774 2862 2811 1 2 ND2 $T=719200 598200 0 0 $X=719200 $Y=597820
X1838 2871 2909 2865 1 2 ND2 $T=726640 557880 1 180 $X=724780 $Y=557500
X1839 2876 395 2860 1 2 ND2 $T=727260 547800 1 0 $X=727260 $Y=542380
X1840 2958 2954 2901 1 2 ND2 $T=733460 588120 1 180 $X=731600 $Y=587740
X1841 2957 2958 2962 1 2 ND2 $T=735320 588120 1 180 $X=733460 $Y=587740
X1842 394 3011 3017 1 2 ND2 $T=739660 688920 1 0 $X=739660 $Y=683500
X1843 3015 3024 2959 1 2 ND2 $T=740900 588120 0 0 $X=740900 $Y=587740
X1844 3018 413 2980 1 2 ND2 $T=747720 547800 1 0 $X=747720 $Y=542380
X1845 415 3094 3080 1 2 ND2 $T=752060 668760 1 180 $X=750200 $Y=668380
X1846 3037 3101 3073 1 2 ND2 $T=755160 547800 1 180 $X=753300 $Y=547420
X1847 2918 3093 3102 1 2 ND2 $T=754540 628440 1 0 $X=754540 $Y=623020
X1848 3112 3110 3094 1 2 ND2 $T=756400 668760 0 180 $X=754540 $Y=663340
X1849 3113 3100 404 1 2 ND2 $T=756400 699000 1 180 $X=754540 $Y=698620
X1850 3062 3111 425 1 2 ND2 $T=758260 678840 0 0 $X=758260 $Y=678460
X1851 2919 3152 3035 1 2 ND2 $T=764460 658680 0 180 $X=762600 $Y=653260
X1852 3105 3185 3060 1 2 ND2 $T=767560 648600 0 180 $X=765700 $Y=643180
X1853 2898 3186 2788 1 2 ND2 $T=767560 658680 1 180 $X=765700 $Y=658300
X1854 2701 3181 3162 1 2 ND2 $T=768800 598200 0 180 $X=766940 $Y=592780
X1855 3222 3208 3189 1 2 ND2 $T=770660 638520 0 180 $X=768800 $Y=633100
X1856 3149 3217 3155 1 2 ND2 $T=770660 648600 0 180 $X=768800 $Y=643180
X1857 3191 3240 3005 1 2 ND2 $T=774380 608280 0 180 $X=772520 $Y=602860
X1858 3198 430 3233 1 2 ND2 $T=776240 547800 0 180 $X=774380 $Y=542380
X1859 3196 3275 3248 1 2 ND2 $T=779960 567960 1 180 $X=778100 $Y=567580
X1860 3257 3284 3302 1 2 ND2 $T=782440 699000 1 0 $X=782440 $Y=693580
X1861 3263 3302 3103 1 2 ND2 $T=784300 699000 1 180 $X=782440 $Y=698620
X1862 3313 3320 3265 1 2 ND2 $T=788640 628440 1 180 $X=786780 $Y=628060
X1863 3255 437 3286 1 2 ND2 $T=789880 547800 1 180 $X=788020 $Y=547420
X1864 3303 3361 3322 1 2 ND2 $T=792360 668760 0 180 $X=790500 $Y=663340
X1865 3329 3360 3336 1 2 ND2 $T=793600 567960 0 180 $X=791740 $Y=562540
X1866 3316 3379 2971 1 2 ND2 $T=795460 598200 0 180 $X=793600 $Y=592780
X1867 3287 3390 3387 1 2 ND2 $T=796700 588120 0 0 $X=796700 $Y=587740
X1868 3342 3394 3378 1 2 ND2 $T=799180 688920 1 180 $X=797320 $Y=688540
X1869 3333 3400 2985 1 2 ND2 $T=801040 638520 0 180 $X=799180 $Y=633100
X1870 3395 3416 3321 1 2 ND2 $T=802280 648600 1 180 $X=800420 $Y=648220
X1871 3310 3419 3325 1 2 ND2 $T=802280 709080 0 180 $X=800420 $Y=703660
X1872 3381 3410 3314 1 2 ND2 $T=801040 557880 1 0 $X=801040 $Y=552460
X1873 3338 3405 3409 1 2 ND2 $T=802900 688920 0 180 $X=801040 $Y=683500
X1874 3393 3432 3374 1 2 ND2 $T=804760 618360 1 180 $X=802900 $Y=617980
X1875 3443 3425 3412 1 2 ND2 $T=805380 598200 0 180 $X=803520 $Y=592780
X1876 3417 3438 3376 1 2 ND2 $T=806620 688920 1 180 $X=804760 $Y=688540
X1877 3414 3435 3310 1 2 ND2 $T=807240 709080 0 180 $X=805380 $Y=703660
X1878 3413 3448 3428 1 2 ND2 $T=807860 699000 0 180 $X=806000 $Y=693580
X1879 3438 3452 3457 1 2 ND2 $T=806620 688920 1 0 $X=806620 $Y=683500
X1880 3432 3453 3459 1 2 ND2 $T=807240 618360 1 0 $X=807240 $Y=612940
X1881 3214 3469 3388 1 2 ND2 $T=809100 638520 0 180 $X=807240 $Y=633100
X1882 3456 3471 3217 1 2 ND2 $T=809720 648600 1 180 $X=807860 $Y=648220
X1883 3437 3472 3441 1 2 ND2 $T=809720 678840 0 180 $X=807860 $Y=673420
X1884 3458 3460 3402 1 2 ND2 $T=810340 567960 1 180 $X=808480 $Y=567580
X1885 3414 3422 3325 1 2 ND2 $T=808480 709080 1 0 $X=808480 $Y=703660
X1886 3476 3488 3477 1 2 ND2 $T=815300 709080 1 180 $X=813440 $Y=708700
X1887 3405 3519 3489 1 2 ND2 $T=817160 678840 0 0 $X=817160 $Y=678460
X1888 3499 3512 3504 1 2 ND2 $T=817780 688920 0 0 $X=817780 $Y=688540
X1889 3497 3543 3448 1 2 ND2 $T=824600 688920 1 180 $X=822740 $Y=688540
X1890 3401 3553 3345 1 2 ND2 $T=826460 668760 1 0 $X=826460 $Y=663340
X1891 2223 3556 466 1 2 ND2 $T=828940 618360 1 180 $X=827080 $Y=617980
X1892 3555 3571 3546 1 2 ND2 $T=832040 618360 0 180 $X=830180 $Y=612940
X1893 3499 3558 3497 1 2 ND2 $T=830800 688920 0 0 $X=830800 $Y=688540
X1894 3545 3579 3571 1 2 ND2 $T=834520 618360 0 180 $X=832660 $Y=612940
X1895 473 3582 471 1 2 ND2 $T=834520 709080 1 180 $X=832660 $Y=708700
X1896 3552 3603 3566 1 2 ND2 $T=835760 608280 0 0 $X=835760 $Y=607900
X1897 3529 3602 3583 1 2 ND2 $T=836380 588120 0 0 $X=836380 $Y=587740
X1898 3604 3601 476 1 2 ND2 $T=838240 709080 0 180 $X=836380 $Y=703660
X1899 3565 3624 3594 1 2 ND2 $T=840720 567960 1 180 $X=838860 $Y=567580
X1900 3610 3625 3603 1 2 ND2 $T=840100 608280 0 0 $X=840100 $Y=607900
X1901 3539 3630 3636 1 2 ND2 $T=841960 598200 1 0 $X=841960 $Y=592780
X1902 486 3646 485 1 2 ND2 $T=845060 557880 0 180 $X=843200 $Y=552460
X1903 3623 3627 3599 1 2 ND2 $T=843200 709080 1 0 $X=843200 $Y=703660
X1904 3622 3638 3617 1 2 ND2 $T=844440 699000 1 0 $X=844440 $Y=693580
X1905 3631 3652 3646 1 2 ND2 $T=845060 557880 0 0 $X=845060 $Y=557500
X1906 3640 3669 3619 1 2 ND2 $T=848160 578040 1 180 $X=846300 $Y=577660
X1907 3666 3672 3630 1 2 ND2 $T=848160 598200 1 0 $X=848160 $Y=592780
X1908 488 3674 480 1 2 ND2 $T=851260 547800 0 180 $X=849400 $Y=542380
X1909 3671 3644 3655 1 2 ND2 $T=851880 699000 1 180 $X=850020 $Y=698620
X1910 3653 3695 3660 1 2 ND2 $T=857460 557880 0 180 $X=855600 $Y=552460
X1911 3693 3697 3624 1 2 ND2 $T=857460 567960 1 180 $X=855600 $Y=567580
X1912 3678 505 3695 1 2 ND2 $T=859320 547800 1 180 $X=857460 $Y=547420
X1913 3739 3745 3710 1 2 ND2 $T=871100 557880 1 180 $X=869240 $Y=557500
X1914 3765 3743 3740 1 2 ND2 $T=872340 578040 1 180 $X=870480 $Y=577660
X1915 3729 3759 3708 1 2 ND2 $T=872340 658680 1 180 $X=870480 $Y=658300
X1916 3776 3738 3769 1 2 ND2 $T=873580 547800 1 0 $X=873580 $Y=542380
X1917 3779 3760 3720 1 2 ND2 $T=875440 567960 1 180 $X=873580 $Y=567580
X1918 3763 3744 3774 1 2 ND2 $T=874200 668760 1 0 $X=874200 $Y=663340
X1919 3785 3766 3798 1 2 ND2 $T=875440 699000 1 0 $X=875440 $Y=693580
X1920 3781 3741 3794 1 2 ND2 $T=876060 658680 1 0 $X=876060 $Y=653260
X1921 3814 3794 3799 1 2 ND2 $T=879780 668760 0 180 $X=877920 $Y=663340
X1922 3785 3824 3749 1 2 ND2 $T=879160 699000 0 0 $X=879160 $Y=698620
X1923 3821 3815 3804 1 2 ND2 $T=881640 567960 1 180 $X=879780 $Y=567580
X1924 3806 3822 3793 1 2 ND2 $T=880400 578040 0 0 $X=880400 $Y=577660
X1925 3746 3833 3811 1 2 ND2 $T=882260 648600 0 180 $X=880400 $Y=643180
X1926 3837 3829 3828 1 2 ND2 $T=884120 638520 0 180 $X=882260 $Y=633100
X1927 3816 3854 3791 1 2 ND2 $T=885980 588120 0 180 $X=884120 $Y=582700
X1928 3835 3841 528 1 2 ND2 $T=884740 567960 1 0 $X=884740 $Y=562540
X1929 3844 3798 3840 1 2 ND2 $T=885980 699000 1 0 $X=885980 $Y=693580
X1930 3850 3826 3839 1 2 ND2 $T=886600 658680 0 0 $X=886600 $Y=658300
X1931 3872 3828 3865 1 2 ND2 $T=890940 658680 1 180 $X=889080 $Y=658300
X1932 3885 3843 3932 1 2 ND2 $T=893420 648600 0 0 $X=893420 $Y=648220
X1933 3906 3901 3846 1 2 ND2 $T=895900 578040 0 180 $X=894040 $Y=572620
X1934 3855 3889 3753 1 2 ND2 $T=894040 588120 0 0 $X=894040 $Y=587740
X1935 3893 3892 3905 1 2 ND2 $T=894040 688920 0 0 $X=894040 $Y=688540
X1936 3892 3912 3881 1 2 ND2 $T=895900 688920 1 0 $X=895900 $Y=683500
X1937 3897 3905 3933 1 2 ND2 $T=896520 699000 1 0 $X=896520 $Y=693580
X1938 535 3949 538 1 2 ND2 $T=897140 709080 0 0 $X=897140 $Y=708700
X1939 538 3942 537 1 2 ND2 $T=899620 719160 0 180 $X=897760 $Y=713740
X1940 3937 3911 3934 1 2 ND2 $T=899620 668760 1 0 $X=899620 $Y=663340
X1941 535 3964 537 1 2 ND2 $T=902720 719160 0 180 $X=900860 $Y=713740
X1942 3959 3948 3967 1 2 ND2 $T=902720 638520 1 0 $X=902720 $Y=633100
X1943 3896 3956 3991 1 2 ND2 $T=903960 588120 0 0 $X=903960 $Y=587740
X1944 3968 3967 3953 1 2 ND2 $T=905200 658680 1 0 $X=905200 $Y=653260
X1945 3985 3977 4003 1 2 ND2 $T=907060 567960 1 0 $X=907060 $Y=562540
X1946 3962 3944 3969 1 2 ND2 $T=909540 699000 0 180 $X=907680 $Y=693580
X1947 4000 3982 4011 1 2 ND2 $T=908920 658680 1 0 $X=908920 $Y=653260
X1948 3979 4007 3831 1 2 ND2 $T=912020 598200 1 180 $X=910160 $Y=597820
X1949 4017 3999 3923 1 2 ND2 $T=912640 567960 0 0 $X=912640 $Y=567580
X1950 4019 3993 4044 1 2 ND2 $T=913260 648600 1 0 $X=913260 $Y=643180
X1951 4043 4026 4024 1 2 ND2 $T=915120 699000 0 180 $X=913260 $Y=693580
X1952 4025 4028 3992 1 2 ND2 $T=913880 557880 0 0 $X=913880 $Y=557500
X1953 3983 4052 4034 1 2 ND2 $T=916980 678840 1 180 $X=915120 $Y=678460
X1954 4057 4044 4036 1 2 ND2 $T=918220 648600 0 0 $X=918220 $Y=648220
X1955 4072 4074 4100 1 2 ND2 $T=921320 648600 1 0 $X=921320 $Y=643180
X1956 4075 4090 4061 1 2 ND2 $T=923800 567960 0 180 $X=921940 $Y=562540
X1957 573 4112 4087 1 2 ND2 $T=925660 547800 1 180 $X=923800 $Y=547420
X1958 4082 4108 3823 1 2 ND2 $T=925660 588120 1 180 $X=923800 $Y=587740
X1959 4037 4100 4084 1 2 ND2 $T=923800 648600 0 0 $X=923800 $Y=648220
X1960 4078 4117 4099 1 2 ND2 $T=926280 598200 0 180 $X=924420 $Y=592780
X1961 4105 4068 4113 1 2 ND2 $T=925040 557880 0 0 $X=925040 $Y=557500
X1962 4116 4126 4105 1 2 ND2 $T=927520 578040 0 180 $X=925660 $Y=572620
X1963 4110 4062 4128 1 2 ND2 $T=926280 648600 1 0 $X=926280 $Y=643180
X1964 4106 4070 4086 1 2 ND2 $T=929380 688920 1 180 $X=927520 $Y=688540
X1965 4136 4131 4116 1 2 ND2 $T=930620 567960 1 180 $X=928760 $Y=567580
X1966 4116 4147 4097 1 2 ND2 $T=930620 578040 1 180 $X=928760 $Y=577660
X1967 4135 4081 4159 1 2 ND2 $T=930620 638520 0 0 $X=930620 $Y=638140
X1968 4151 4125 4145 1 2 ND2 $T=934340 648600 1 0 $X=934340 $Y=643180
X1969 577 4156 576 1 2 ND2 $T=936200 699000 1 180 $X=934340 $Y=698620
X1970 4152 4172 4156 1 2 ND2 $T=938060 699000 0 180 $X=936200 $Y=693580
X1971 4172 4171 4154 1 2 ND2 $T=938680 699000 1 180 $X=936820 $Y=698620
X1972 4150 4144 4174 1 2 ND2 $T=938060 628440 0 0 $X=938060 $Y=628060
X1973 4175 4174 4166 1 2 ND2 $T=939920 648600 1 0 $X=939920 $Y=643180
X1974 4191 4184 4199 1 2 ND2 $T=944260 638520 0 0 $X=944260 $Y=638140
X1975 4183 4211 4201 1 2 ND2 $T=949840 699000 1 180 $X=947980 $Y=698620
X1976 4222 4214 4234 1 2 ND2 $T=952320 678840 1 0 $X=952320 $Y=673420
X1977 4226 4234 602 1 2 ND2 $T=953560 709080 1 0 $X=953560 $Y=703660
X1978 4129 4253 4237 1 2 ND2 $T=959760 678840 1 180 $X=957900 $Y=678460
X1979 604 4250 607 1 2 ND2 $T=958520 719160 1 0 $X=958520 $Y=713740
X1980 609 4257 611 1 2 ND2 $T=967820 709080 1 0 $X=967820 $Y=703660
X1981 4264 4332 4300 1 2 ND2 $T=981460 688920 0 180 $X=979600 $Y=683500
X1982 702 727 1 741 2 743 OAI12HS $T=279620 638520 0 180 $X=275900 $Y=633100
X1983 782 772 1 805 2 798 OAI12HS $T=290780 598200 1 0 $X=290780 $Y=592780
X1984 825 818 1 806 2 778 OAI12HS $T=296360 648600 1 180 $X=292640 $Y=648220
X1985 827 823 1 792 2 806 OAI12HS $T=298220 658680 1 0 $X=298220 $Y=653260
X1986 912 900 1 915 2 21 OAI12HS $T=313100 547800 0 0 $X=313100 $Y=547420
X1987 944 938 1 928 2 926 OAI12HS $T=318680 608280 0 180 $X=314960 $Y=602860
X1988 918 945 1 935 2 904 OAI12HS $T=320540 638520 1 180 $X=316820 $Y=638140
X1989 947 952 1 933 2 25 OAI12HS $T=318680 547800 1 0 $X=318680 $Y=542380
X1990 965 952 1 956 2 975 OAI12HS $T=322400 547800 0 0 $X=322400 $Y=547420
X1991 923 28 1 912 2 969 OAI12HS $T=326120 557880 1 0 $X=326120 $Y=552460
X1992 918 1017 1 970 2 1010 OAI12HS $T=334800 628440 1 180 $X=331080 $Y=628060
X1993 31 34 1 1003 2 32 OAI12HS $T=335420 547800 0 180 $X=331700 $Y=542380
X1994 1101 1094 1 1088 2 1042 OAI12HS $T=347200 608280 0 180 $X=343480 $Y=602860
X1995 1114 954 1 979 2 1120 OAI12HS $T=353400 567960 0 180 $X=349680 $Y=562540
X1996 1111 1117 1 1137 2 1088 OAI12HS $T=350920 608280 1 0 $X=350920 $Y=602860
X1997 1132 1044 1 1031 2 1156 OAI12HS $T=358360 557880 1 180 $X=354640 $Y=557500
X1998 1180 867 1 983 2 1064 OAI12HS $T=358980 618360 1 180 $X=355260 $Y=617980
X1999 1171 1167 1 1142 2 1151 OAI12HS $T=361460 557880 0 180 $X=357740 $Y=552460
X2000 1085 1162 1 1114 2 1178 OAI12HS $T=357740 567960 0 0 $X=357740 $Y=567580
X2001 1224 1233 1 1246 2 1197 OAI12HS $T=368280 588120 0 0 $X=368280 $Y=587740
X2002 1220 61 1 1167 2 1284 OAI12HS $T=373860 547800 0 0 $X=373860 $Y=547420
X2003 1270 1273 1 1237 2 1289 OAI12HS $T=374480 567960 0 0 $X=374480 $Y=567580
X2004 1272 1273 1 1254 2 1292 OAI12HS $T=375100 567960 1 0 $X=375100 $Y=562540
X2005 1219 1263 1 1290 2 1246 OAI12HS $T=376340 588120 0 0 $X=376340 $Y=587740
X2006 1285 1273 1 1232 2 1307 OAI12HS $T=376960 557880 0 0 $X=376960 $Y=557500
X2007 1325 1319 1 1310 2 62 OAI12HS $T=385020 547800 0 180 $X=381300 $Y=542380
X2008 1336 61 1 1325 2 1377 OAI12HS $T=391840 547800 1 0 $X=391840 $Y=542380
X2009 1386 1393 1 1403 2 1334 OAI12HS $T=396800 699000 0 0 $X=396800 $Y=698620
X2010 1335 1395 1 1385 2 1387 OAI12HS $T=400520 709080 1 180 $X=396800 $Y=708700
X2011 1240 1312 1 1399 2 1398 OAI12HS $T=397420 638520 0 0 $X=397420 $Y=638140
X2012 1387 78 1 80 2 1403 OAI12HS $T=400520 709080 1 0 $X=400520 $Y=703660
X2013 1414 1419 1 1424 2 79 OAI12HS $T=401760 547800 1 0 $X=401760 $Y=542380
X2014 1446 1419 1 1464 2 95 OAI12HS $T=409820 547800 1 0 $X=409820 $Y=542380
X2015 1394 1395 1 1463 2 1469 OAI12HS $T=409820 709080 0 0 $X=409820 $Y=708700
X2016 1517 99 1 1501 2 1482 OAI12HS $T=422840 547800 1 180 $X=419120 $Y=547420
X2017 1718 1686 1 1705 2 1709 OAI12HS $T=465620 557880 0 180 $X=461900 $Y=552460
X2018 1748 1713 1 1710 2 1738 OAI12HS $T=470580 578040 0 180 $X=466860 $Y=572620
X2019 1756 1746 1 1737 2 1145 OAI12HS $T=471820 557880 0 180 $X=468100 $Y=552460
X2020 1731 1759 1 1718 2 1753 OAI12HS $T=473060 557880 1 180 $X=469340 $Y=557500
X2021 1758 1749 1 1715 2 1767 OAI12HS $T=471820 618360 1 0 $X=471820 $Y=612940
X2022 1775 1777 1 1766 2 1768 OAI12HS $T=476160 588120 0 180 $X=472440 $Y=582700
X2023 1786 1781 1 1754 2 1774 OAI12HS $T=476780 598200 1 180 $X=473060 $Y=597820
X2024 1743 1784 1 1775 2 1831 OAI12HS $T=479880 588120 0 0 $X=479880 $Y=587740
X2025 1787 1797 1 1850 2 1810 OAI12HS $T=484840 648600 1 0 $X=484840 $Y=643180
X2026 2165 249 1 2151 2 2157 OAI12HS $T=563580 628440 1 180 $X=559860 $Y=628060
X2027 2767 2789 1 2801 2 2812 OAI12HS $T=710520 699000 0 0 $X=710520 $Y=698620
X2028 2850 2821 1 2804 2 2810 OAI12HS $T=719200 598200 1 180 $X=715480 $Y=597820
X2029 2823 2828 1 2888 2 2902 OAI12HS $T=721680 658680 0 0 $X=721680 $Y=658300
X2030 2863 2892 1 2902 2 2898 OAI12HS $T=723540 668760 1 0 $X=723540 $Y=663340
X2031 2861 2855 1 2820 2 2905 OAI12HS $T=725400 567960 0 0 $X=725400 $Y=567580
X2032 398 394 1 2900 2 2725 OAI12HS $T=729120 709080 0 180 $X=725400 $Y=703660
X2033 2924 2916 1 2894 2 2908 OAI12HS $T=729740 547800 1 180 $X=726020 $Y=547420
X2034 2683 2918 1 2837 2 2891 OAI12HS $T=726020 608280 0 0 $X=726020 $Y=607900
X2035 2939 2946 1 2926 2 2888 OAI12HS $T=730360 658680 1 180 $X=726640 $Y=658300
X2036 2920 384 1 2933 2 2928 OAI12HS $T=727260 678840 1 0 $X=727260 $Y=673420
X2037 2951 2952 1 2928 2 2926 OAI12HS $T=732220 668760 0 180 $X=728500 $Y=663340
X2038 2973 396 1 2903 2 2933 OAI12HS $T=734700 678840 0 180 $X=730980 $Y=673420
X2039 2976 2927 1 2963 2 2978 OAI12HS $T=734700 598200 1 0 $X=734700 $Y=592780
X2040 406 2994 1 367 2 2951 OAI12HS $T=736560 719160 1 0 $X=736560 $Y=713740
X2041 3003 2890 1 2998 2 3028 OAI12HS $T=745240 557880 0 180 $X=741520 $Y=552460
X2042 2927 3040 1 3024 2 3052 OAI12HS $T=743380 588120 0 0 $X=743380 $Y=587740
X2043 3023 3049 1 3028 2 414 OAI12HS $T=745240 547800 0 0 $X=745240 $Y=547420
X2044 3033 3014 1 3011 2 3047 OAI12HS $T=745240 678840 0 0 $X=745240 $Y=678460
X2045 3053 3061 1 3071 2 3079 OAI12HS $T=746480 658680 1 0 $X=746480 $Y=653260
X2046 2937 2955 1 3093 2 3085 OAI12HS $T=750200 628440 0 0 $X=750200 $Y=628060
X2047 3072 3014 1 3100 2 3103 OAI12HS $T=750820 699000 0 0 $X=750820 $Y=698620
X2048 3082 416 1 3101 2 423 OAI12HS $T=751440 547800 1 0 $X=751440 $Y=542380
X2049 3080 415 1 2904 2 3112 OAI12HS $T=752680 668760 0 0 $X=752680 $Y=668380
X2050 2913 3048 1 3110 2 3071 OAI12HS $T=753300 658680 1 0 $X=753300 $Y=653260
X2051 419 412 1 3111 2 3080 OAI12HS $T=753300 678840 0 0 $X=753300 $Y=678460
X2052 3166 2822 1 3076 2 3190 OAI12HS $T=770040 628440 0 180 $X=766320 $Y=623020
X2053 3085 3179 1 3231 2 3222 OAI12HS $T=771280 638520 1 0 $X=771280 $Y=633100
X2054 2785 3226 1 3190 2 3231 OAI12HS $T=771900 628440 1 0 $X=771900 $Y=623020
X2055 3088 3219 1 3215 2 3250 OAI12HS $T=778720 688920 0 180 $X=775000 $Y=683500
X2056 3274 3267 1 3250 2 3253 OAI12HS $T=781200 678840 1 180 $X=777480 $Y=678460
X2057 3103 3263 1 3210 2 3257 OAI12HS $T=781820 699000 1 180 $X=778100 $Y=698620
X2058 3249 3268 1 3275 2 3283 OAI12HS $T=778720 567960 1 0 $X=778720 $Y=562540
X2059 3147 3273 1 3204 2 3313 OAI12HS $T=781820 628440 0 0 $X=781820 $Y=628060
X2060 3298 3312 1 3319 2 3332 OAI12HS $T=785540 588120 1 0 $X=785540 $Y=582700
X2061 3266 3091 1 3320 2 3330 OAI12HS $T=791120 638520 0 180 $X=787400 $Y=633100
X2062 2971 3316 1 3323 2 3318 OAI12HS $T=791740 598200 0 180 $X=788020 $Y=592780
X2063 3344 3353 1 3362 2 3369 OAI12HS $T=791740 709080 0 0 $X=791740 $Y=708700
X2064 3345 3334 1 3361 2 3371 OAI12HS $T=797320 668760 0 180 $X=793600 $Y=663340
X2065 3259 3001 1 441 2 3362 OAI12HS $T=794220 719160 1 0 $X=794220 $Y=713740
X2066 3350 3372 1 3330 2 3388 OAI12HS $T=794840 638520 1 0 $X=794840 $Y=633100
X2067 3364 3384 1 3394 2 3409 OAI12HS $T=796700 688920 1 0 $X=796700 $Y=683500
X2068 3415 3412 1 3432 2 3420 OAI12HS $T=802280 618360 1 0 $X=802280 $Y=612940
X2069 3495 3481 1 3484 2 3526 OAI12HS $T=815920 648600 1 0 $X=815920 $Y=643180
X2070 3606 3542 1 3556 2 3598 OAI12HS $T=839480 618360 1 180 $X=835760 $Y=617980
X2071 3582 3596 1 3601 2 3605 OAI12HS $T=835760 699000 0 0 $X=835760 $Y=698620
X2072 3612 3609 1 3603 2 3621 OAI12HS $T=845680 608280 0 180 $X=841960 $Y=602860
X2073 3627 3635 1 3644 2 3629 OAI12HS $T=842580 699000 0 0 $X=842580 $Y=698620
X2074 3650 3643 1 3627 2 3642 OAI12HS $T=846920 678840 1 180 $X=843200 $Y=678460
X2075 3638 479 1 3639 2 3663 OAI12HS $T=843820 688920 0 0 $X=843820 $Y=688540
X2076 3630 3589 1 3602 2 3647 OAI12HS $T=848160 588120 1 180 $X=844440 $Y=587740
X2077 3646 3667 1 3674 2 3670 OAI12HS $T=848160 547800 0 0 $X=848160 $Y=547420
X2078 3626 3668 1 3646 2 3664 OAI12HS $T=851880 557880 1 180 $X=848160 $Y=557500
X2079 3669 3651 1 3624 2 3645 OAI12HS $T=848780 567960 0 0 $X=848780 $Y=567580
X2080 3738 511 1 3756 2 512 OAI12HS $T=868000 547800 1 0 $X=868000 $Y=542380
X2081 3760 3751 1 3743 2 3750 OAI12HS $T=871720 567960 0 180 $X=868000 $Y=562540
X2082 3731 3757 1 3759 2 3724 OAI12HS $T=869860 638520 0 0 $X=869860 $Y=638140
X2083 516 3730 1 3745 2 3768 OAI12HS $T=874200 547800 1 180 $X=870480 $Y=547420
X2084 3754 3757 1 3770 2 3733 OAI12HS $T=871720 648600 1 0 $X=871720 $Y=643180
X2085 3759 3762 1 3744 2 3773 OAI12HS $T=871720 658680 1 0 $X=871720 $Y=653260
X2086 3780 3786 1 3789 2 3787 OAI12HS $T=874820 638520 0 0 $X=874820 $Y=638140
X2087 3784 3801 1 3760 2 3813 OAI12HS $T=877300 557880 0 0 $X=877300 $Y=557500
X2088 3833 3786 1 3809 2 3807 OAI12HS $T=882880 638520 1 180 $X=879160 $Y=638140
X2089 3794 3819 1 3826 2 3818 OAI12HS $T=879780 658680 1 0 $X=879780 $Y=653260
X2090 3812 509 1 3803 2 3827 OAI12HS $T=885980 547800 0 180 $X=882260 $Y=542380
X2091 3805 509 1 3825 2 3879 OAI12HS $T=882260 557880 1 0 $X=882260 $Y=552460
X2092 3860 3786 1 3847 2 3853 OAI12HS $T=888460 638520 0 180 $X=884740 $Y=633100
X2093 3822 3832 1 3854 2 3868 OAI12HS $T=886600 578040 0 0 $X=886600 $Y=577660
X2094 3843 3809 1 3880 2 3861 OAI12HS $T=889080 648600 0 0 $X=889080 $Y=648220
X2095 541 534 1 3876 2 3897 OAI12HS $T=895900 699000 1 180 $X=892180 $Y=698620
X2096 3877 3926 1 3841 2 3902 OAI12HS $T=897140 567960 0 180 $X=893420 $Y=562540
X2097 3899 3786 1 3913 2 3918 OAI12HS $T=894040 638520 1 0 $X=894040 $Y=633100
X2098 3900 3786 1 3914 2 3931 OAI12HS $T=894040 638520 0 0 $X=894040 $Y=638140
X2099 3828 3910 1 3911 2 3909 OAI12HS $T=894660 658680 1 0 $X=894660 $Y=653260
X2100 3916 3929 1 3938 2 3888 OAI12HS $T=897140 588120 1 0 $X=897140 $Y=582700
X2101 3935 3929 1 3943 2 3965 OAI12HS $T=900860 567960 0 0 $X=900860 $Y=567580
X2102 3952 3958 1 3967 2 3947 OAI12HS $T=901480 648600 1 0 $X=901480 $Y=643180
X2103 3967 3975 1 3982 2 3941 OAI12HS $T=904580 648600 0 0 $X=904580 $Y=648220
X2104 3977 3981 1 3989 2 555 OAI12HS $T=905820 557880 0 0 $X=905820 $Y=557500
X2105 4001 3864 1 3976 2 3987 OAI12HS $T=909540 638520 1 180 $X=905820 $Y=638140
X2106 3972 3981 1 3999 2 3990 OAI12HS $T=907060 578040 1 0 $X=907060 $Y=572620
X2107 3980 3984 1 3997 2 3969 OAI12HS $T=907060 699000 0 0 $X=907060 $Y=698620
X2108 549 3963 1 3925 2 3997 OAI12HS $T=907680 709080 1 0 $X=907680 $Y=703660
X2109 3901 3929 1 3908 2 4033 OAI12HS $T=918840 578040 0 180 $X=915120 $Y=572620
X2110 4051 566 1 4050 2 4077 OAI12HS $T=923800 709080 0 180 $X=920080 $Y=703660
X2111 4068 3908 1 4088 2 4059 OAI12HS $T=920700 557880 0 0 $X=920700 $Y=557500
X2112 4083 4022 1 4062 2 4098 OAI12HS $T=922560 628440 0 0 $X=922560 $Y=628060
X2113 4081 4022 1 4095 2 4069 OAI12HS $T=922560 638520 1 0 $X=922560 $Y=633100
X2114 4064 4095 1 4100 2 4018 OAI12HS $T=922560 638520 0 0 $X=922560 $Y=638140
X2115 4109 4066 1 4077 2 4086 OAI12HS $T=926280 699000 1 180 $X=922560 $Y=698620
X2116 4046 4120 1 4090 2 4111 OAI12HS $T=930000 567960 0 180 $X=926280 $Y=562540
X2117 4134 4022 1 4115 2 4122 OAI12HS $T=930000 628440 0 180 $X=926280 $Y=623020
X2118 4062 4118 1 4125 2 4124 OAI12HS $T=926280 638520 0 0 $X=926280 $Y=638140
X2119 4108 4127 1 4117 2 4119 OAI12HS $T=927520 588120 0 0 $X=927520 $Y=587740
X2120 4126 3929 1 4139 2 4091 OAI12HS $T=928140 578040 1 0 $X=928140 $Y=572620
X2121 4090 4130 1 4112 2 4138 OAI12HS $T=930000 557880 1 0 $X=930000 $Y=552460
X2122 4131 3929 1 4148 2 4142 OAI12HS $T=930000 567960 1 0 $X=930000 $Y=562540
X2123 4141 4022 1 4149 2 4163 OAI12HS $T=930620 628440 1 0 $X=930620 $Y=623020
X2124 576 577 1 4085 2 4152 OAI12HS $T=930620 699000 0 0 $X=930620 $Y=698620
X2125 4147 3929 1 4123 2 4158 OAI12HS $T=931860 578040 0 0 $X=931860 $Y=577660
X2126 4174 4177 1 4184 2 4161 OAI12HS $T=939920 638520 0 0 $X=939920 $Y=638140
X2127 4242 4243 1 4228 2 606 OAI12HS $T=957280 547800 0 0 $X=957280 $Y=547420
X2128 4271 4260 1 4275 2 610 OAI12HS $T=964720 547800 1 0 $X=964720 $Y=542380
X2129 686 678 1 677 2 NR2T $T=259780 628440 1 180 $X=254820 $Y=628060
X2130 767 762 1 771 2 NR2T $T=287680 618360 0 180 $X=282720 $Y=612940
X2131 813 775 1 784 2 NR2T $T=295120 668760 0 180 $X=290160 $Y=663340
X2132 809 813 1 847 2 NR2T $T=295740 608280 1 0 $X=295740 $Y=602860
X2133 916 966 1 960 2 NR2T $T=323020 588120 0 180 $X=318060 $Y=582700
X2134 960 941 1 967 2 NR2T $T=324260 588120 1 180 $X=319300 $Y=587740
X2135 1039 1079 1 42 2 NR2T $T=339760 709080 0 0 $X=339760 $Y=708700
X2136 1128 1129 1 1122 2 NR2T $T=352780 588120 1 180 $X=347820 $Y=587740
X2137 959 1128 1 1125 2 NR2T $T=353400 578040 1 180 $X=348440 $Y=577660
X2138 1079 48 1 1107 2 NR2T $T=350300 709080 0 0 $X=350300 $Y=708700
X2139 1062 1141 1 1154 2 NR2T $T=357740 699000 1 180 $X=352780 $Y=698620
X2140 3315 3328 1 3278 2 NR2T $T=790500 547800 0 180 $X=785540 $Y=542380
X2141 3431 3295 1 3383 2 NR2T $T=801040 608280 1 180 $X=796080 $Y=607900
X2142 3450 3436 1 3424 2 NR2T $T=807860 588120 1 0 $X=807860 $Y=582700
X2143 3480 3436 1 3424 2 NR2T $T=813440 578040 0 0 $X=813440 $Y=577660
X2144 3530 3506 1 3449 2 NR2T $T=822120 618360 1 0 $X=822120 $Y=612940
X2145 4307 4338 1 621 2 NR2T $T=983320 719160 1 0 $X=983320 $Y=713740
X2146 4338 4312 1 4329 2 NR2T $T=984560 709080 1 0 $X=984560 $Y=703660
X2147 710 1 715 703 2 720 ND3 $T=267840 578040 0 0 $X=267840 $Y=577660
X2148 739 1 756 764 2 748 ND3 $T=280240 578040 1 0 $X=280240 $Y=572620
X2149 790 1 793 784 2 812 ND3 $T=290160 688920 1 0 $X=290160 $Y=683500
X2150 1027 1 1005 1004 2 1007 ND3 $T=329220 578040 0 0 $X=329220 $Y=577660
X2151 991 1 1035 1027 2 959 ND3 $T=336040 578040 1 180 $X=333560 $Y=577660
X2152 1112 1 1099 1093 2 1062 ND3 $T=347820 699000 1 180 $X=345340 $Y=698620
X2153 1093 1 1100 1078 2 46 ND3 $T=345960 709080 1 0 $X=345960 $Y=703660
X2154 115 1 122 1650 2 125 ND3 $T=449500 719160 1 0 $X=449500 $Y=713740
X2155 2909 1 2917 393 2 2889 ND3 $T=726020 557880 1 0 $X=726020 $Y=552460
X2156 3402 1 3423 3380 2 3407 ND3 $T=803520 567960 1 180 $X=801040 $Y=567580
X2157 3419 1 3422 3428 2 3435 ND3 $T=802900 709080 1 0 $X=802900 $Y=703660
X2158 3443 1 3450 3426 2 3454 ND3 $T=806620 598200 1 0 $X=806620 $Y=592780
X2159 3458 1 3486 3407 2 3454 ND3 $T=814060 567960 1 180 $X=811580 $Y=567580
X2160 3462 1 3480 3483 2 3454 ND3 $T=811580 598200 1 0 $X=811580 $Y=592780
X2161 3497 1 3505 3541 2 3544 ND3 $T=824600 699000 1 0 $X=824600 $Y=693580
X2162 3541 1 3448 3549 2 3558 ND3 $T=826460 688920 0 0 $X=826460 $Y=688540
X2163 3698 1 3699 3714 2 3696 ND3 $T=856840 588120 0 0 $X=856840 $Y=587740
X2164 3942 1 3949 3963 2 3964 ND3 $T=900240 709080 0 0 $X=900240 $Y=708700
X2165 4034 1 3862 4015 2 3970 ND3 $T=911400 678840 1 180 $X=908920 $Y=678460
X2166 4052 1 4015 4067 2 4026 ND3 $T=917600 678840 0 0 $X=917600 $Y=678460
X2167 4234 1 4241 4254 2 4253 ND3 $T=957280 678840 1 0 $X=957280 $Y=673420
X2168 611 1 4274 4289 2 4279 ND3 $T=966580 678840 0 0 $X=966580 $Y=678460
X2169 609 1 4249 4279 2 4162 ND3 $T=967200 688920 1 0 $X=967200 $Y=683500
X2170 4314 1 4249 4310 2 4162 ND3 $T=974020 688920 0 0 $X=974020 $Y=688540
X2171 4340 1 4332 4311 2 4293 ND3 $T=983320 688920 1 0 $X=983320 $Y=683500
X2172 4312 1 4334 4347 2 4310 ND3 $T=984560 688920 0 0 $X=984560 $Y=688540
X2173 688 712 699 2 1 XNR2HS $T=269700 608280 1 180 $X=264120 $Y=607900
X2174 733 736 737 2 1 XNR2HS $T=273420 618360 1 0 $X=273420 $Y=612940
X2175 723 745 731 2 1 XNR2HS $T=279620 658680 1 180 $X=274040 $Y=658300
X2176 751 746 736 2 1 XNR2HS $T=280240 618360 1 180 $X=274660 $Y=617980
X2177 689 687 745 2 1 XNR2HS $T=285820 658680 1 180 $X=280240 $Y=658300
X2178 778 773 682 2 1 XNR2HS $T=288920 648600 1 180 $X=283340 $Y=648220
X2179 789 774 765 2 1 XNR2HS $T=291400 678840 0 180 $X=285820 $Y=673420
X2180 792 788 689 2 1 XNR2HS $T=292020 658680 1 180 $X=286440 $Y=658300
X2181 827 823 788 2 1 XNR2HS $T=297600 658680 1 180 $X=292020 $Y=658300
X2182 820 845 802 2 1 XNR2HS $T=302560 678840 1 180 $X=296980 $Y=678460
X2183 854 829 846 2 1 XNR2HS $T=304420 688920 1 180 $X=298840 $Y=688540
X2184 855 811 858 2 1 XNR2HS $T=301940 588120 0 0 $X=301940 $Y=587740
X2185 877 902 854 2 1 XNR2HS $T=311860 688920 0 180 $X=306280 $Y=683500
X2186 871 914 861 2 1 XNR2HS $T=314340 668760 1 180 $X=308760 $Y=668380
X2187 932 871 864 2 1 XNR2HS $T=316820 668760 0 180 $X=311240 $Y=663340
X2188 888 907 902 2 1 XNR2HS $T=311860 678840 0 0 $X=311860 $Y=678460
X2189 939 914 844 2 1 XNR2HS $T=318680 658680 0 180 $X=313100 $Y=653260
X2190 944 938 925 2 1 XNR2HS $T=319300 598200 1 180 $X=313720 $Y=597820
X2191 925 928 941 2 1 XNR2HS $T=314340 598200 1 0 $X=314340 $Y=592780
X2192 964 958 839 2 1 XNR2HS $T=322400 688920 0 180 $X=316820 $Y=683500
X2193 974 976 872 2 1 XNR2HS $T=325500 648600 1 180 $X=319920 $Y=648220
X2194 957 969 978 2 1 XNR2HS $T=320540 557880 1 0 $X=320540 $Y=552460
X2195 903 975 980 2 1 XNR2HS $T=322400 547800 1 0 $X=322400 $Y=542380
X2196 939 1001 945 2 1 XNR2HS $T=331080 658680 1 180 $X=325500 $Y=658300
X2197 998 994 944 2 1 XNR2HS $T=332940 678840 0 180 $X=327360 $Y=673420
X2198 997 932 1011 2 1 XNR2HS $T=327980 648600 1 0 $X=327980 $Y=643180
X2199 989 976 875 2 1 XNR2HS $T=333560 658680 0 180 $X=327980 $Y=653260
X2200 999 1004 1014 2 1 XNR2HS $T=328600 578040 1 0 $X=328600 $Y=572620
X2201 1000 996 1015 2 1 XNR2HS $T=328600 598200 0 0 $X=328600 $Y=597820
X2202 1025 871 962 2 1 XNR2HS $T=334800 668760 1 180 $X=329220 $Y=668380
X2203 997 914 1021 2 1 XNR2HS $T=329840 648600 0 0 $X=329840 $Y=648220
X2204 977 997 1037 2 1 XNR2HS $T=343480 648600 1 180 $X=337900 $Y=648220
X2205 1001 1018 984 2 1 XNR2HS $T=338520 658680 0 0 $X=338520 $Y=658300
X2206 1080 1078 1068 2 1 XNR2HS $T=344720 709080 0 180 $X=339140 $Y=703660
X2207 1070 1072 1082 2 1 XNR2HS $T=340380 608280 0 0 $X=340380 $Y=607900
X2208 997 989 1051 2 1 XNR2HS $T=345960 638520 0 180 $X=340380 $Y=633100
X2209 1073 1089 1070 2 1 XNR2HS $T=346580 618360 1 180 $X=341000 $Y=617980
X2210 1095 1091 1073 2 1 XNR2HS $T=346580 638520 1 180 $X=341000 $Y=638140
X2211 1092 963 1066 2 1 XNR2HS $T=347820 658680 0 0 $X=347820 $Y=658300
X2212 50 1092 1050 2 1 XNR2HS $T=353400 678840 1 180 $X=347820 $Y=678460
X2213 1137 1138 1115 2 1 XNR2HS $T=355260 598200 1 180 $X=349680 $Y=597820
X2214 1111 1117 1138 2 1 XNR2HS $T=349680 608280 0 0 $X=349680 $Y=607900
X2215 1147 974 1059 2 1 XNR2HS $T=355880 648600 0 180 $X=350300 $Y=643180
X2216 1092 1131 1104 2 1 XNR2HS $T=357120 658680 0 180 $X=351540 $Y=653260
X2217 1092 1155 1086 2 1 XNR2HS $T=357740 668760 0 180 $X=352160 $Y=663340
X2218 1150 1139 1102 2 1 XNR2HS $T=358360 628440 1 180 $X=352780 $Y=628060
X2219 1148 1159 1168 2 1 XNR2HS $T=355880 578040 1 0 $X=355880 $Y=572620
X2220 1179 983 1097 2 1 XNR2HS $T=362700 628440 0 180 $X=357120 $Y=623020
X2221 1204 1214 1198 2 1 XNR2HS $T=367660 688920 1 180 $X=362080 $Y=688540
X2222 1147 1223 1164 2 1 XNR2HS $T=368900 638520 1 180 $X=363320 $Y=638140
X2223 1109 1018 1221 2 1 XNR2HS $T=363320 658680 1 0 $X=363320 $Y=653260
X2224 1169 1206 1203 2 1 XNR2HS $T=363940 598200 0 0 $X=363940 $Y=597820
X2225 1195 1227 1205 2 1 XNR2HS $T=370140 608280 1 180 $X=364560 $Y=607900
X2226 1213 971 1238 2 1 XNR2HS $T=366420 578040 0 0 $X=366420 $Y=577660
X2227 1263 1219 1239 2 1 XNR2HS $T=374480 588120 0 180 $X=368900 $Y=582700
X2228 1259 1230 1263 2 1 XNR2HS $T=375100 608280 1 0 $X=375100 $Y=602860
X2229 1018 1155 1252 2 1 XNR2HS $T=380680 658680 0 180 $X=375100 $Y=653260
X2230 1282 1099 1286 2 1 XNR2HS $T=375720 688920 1 0 $X=375720 $Y=683500
X2231 1278 1284 1304 2 1 XNR2HS $T=376960 557880 1 0 $X=376960 $Y=552460
X2232 1105 1289 1308 2 1 XNR2HS $T=377580 578040 1 0 $X=377580 $Y=572620
X2233 1271 1266 1314 2 1 XNR2HS $T=378820 608280 0 0 $X=378820 $Y=607900
X2234 1193 1292 1320 2 1 XNR2HS $T=379440 567960 1 0 $X=379440 $Y=562540
X2235 1207 1307 1328 2 1 XNR2HS $T=381920 557880 0 0 $X=381920 $Y=557500
X2236 1121 1315 1294 2 1 XNR2HS $T=388740 638520 1 180 $X=383160 $Y=638140
X2237 1121 1339 1248 2 1 XNR2HS $T=389360 628440 0 180 $X=383780 $Y=623020
X2238 1342 1356 1348 2 1 XNR2HS $T=393080 598200 1 180 $X=387500 $Y=597820
X2239 1344 1131 1312 2 1 XNR2HS $T=387500 648600 1 0 $X=387500 $Y=643180
X2240 73 67 1340 2 1 XNR2HS $T=393080 709080 1 180 $X=387500 $Y=708700
X2241 1351 1330 1364 2 1 XNR2HS $T=388740 699000 1 0 $X=388740 $Y=693580
X2242 1340 1334 1351 2 1 XNR2HS $T=394940 688920 1 180 $X=389360 $Y=688540
X2243 1378 1371 1247 2 1 XNR2HS $T=394320 618360 0 0 $X=394320 $Y=617980
X2244 1376 1380 1330 2 1 XNR2HS $T=394320 699000 1 0 $X=394320 $Y=693580
X2245 1350 1377 76 2 1 XNR2HS $T=395560 547800 1 0 $X=395560 $Y=542380
X2246 1330 1351 1409 2 1 XNR2HS $T=398660 688920 0 0 $X=398660 $Y=688540
X2247 1372 1398 1423 2 1 XNR2HS $T=399900 638520 1 0 $X=399900 $Y=633100
X2248 1408 1339 1432 2 1 XNR2HS $T=403000 618360 0 0 $X=403000 $Y=617980
X2249 88 85 1395 2 1 XNR2HS $T=409820 709080 1 180 $X=404240 $Y=708700
X2250 1387 78 1445 2 1 XNR2HS $T=404860 709080 1 0 $X=404860 $Y=703660
X2251 1440 1404 1460 2 1 XNR2HS $T=407960 608280 1 0 $X=407960 $Y=602860
X2252 1339 1344 1473 2 1 XNR2HS $T=410440 628440 0 0 $X=410440 $Y=628060
X2253 91 83 1438 2 1 XNR2HS $T=411060 699000 0 0 $X=411060 $Y=698620
X2254 80 1445 1465 2 1 XNR2HS $T=411060 709080 1 0 $X=411060 $Y=703660
X2255 1189 1408 1461 2 1 XNR2HS $T=417260 628440 0 180 $X=411680 $Y=623020
X2256 1438 1442 1476 2 1 XNR2HS $T=420360 688920 1 180 $X=414780 $Y=688540
X2257 1469 100 1507 2 1 XNR2HS $T=417260 699000 0 0 $X=417260 $Y=698620
X2258 1484 1439 1519 2 1 XNR2HS $T=419740 638520 1 0 $X=419740 $Y=633100
X2259 1189 1382 1541 2 1 XNR2HS $T=425320 638520 0 0 $X=425320 $Y=638140
X2260 1378 1536 1540 2 1 XNR2HS $T=427800 628440 1 0 $X=427800 $Y=623020
X2261 1567 1532 1547 2 1 XNR2HS $T=434620 688920 1 180 $X=429040 $Y=688540
X2262 1523 108 1394 2 1 XNR2HS $T=429660 709080 1 0 $X=429660 $Y=703660
X2263 1561 1550 1579 2 1 XNR2HS $T=433380 628440 1 0 $X=433380 $Y=623020
X2264 1573 1570 1591 2 1 XNR2HS $T=434620 598200 1 0 $X=434620 $Y=592780
X2265 118 1598 1583 2 1 XNR2HS $T=440820 699000 1 180 $X=435240 $Y=698620
X2266 1623 1595 1634 2 1 XNR2HS $T=443300 668760 0 0 $X=443300 $Y=668380
X2267 1580 1607 1611 2 1 XNR2HS $T=443300 699000 1 0 $X=443300 $Y=693580
X2268 1610 1655 1652 2 1 XNR2HS $T=452600 618360 0 0 $X=452600 $Y=617980
X2269 131 1667 1678 2 1 XNR2HS $T=455080 709080 0 0 $X=455080 $Y=708700
X2270 1690 1700 1687 2 1 XNR2HS $T=463140 699000 0 180 $X=457560 $Y=693580
X2271 1776 1789 1815 2 1 XNR2HS $T=478020 618360 1 0 $X=478020 $Y=612940
X2272 1806 1783 1830 2 1 XNR2HS $T=480500 567960 0 0 $X=480500 $Y=567580
X2273 1767 1814 1845 2 1 XNR2HS $T=482360 608280 0 0 $X=482360 $Y=607900
X2274 1819 1831 1848 2 1 XNR2HS $T=482980 588120 1 0 $X=482980 $Y=582700
X2275 2626 2640 2647 2 1 XNR2HS $T=683240 588120 0 0 $X=683240 $Y=587740
X2276 2604 2663 2683 2 1 XNR2HS $T=690060 608280 0 0 $X=690060 $Y=607900
X2277 2717 2706 2691 2 1 XNR2HS $T=701220 557880 0 180 $X=695640 $Y=552460
X2278 2642 2631 2709 2 1 XNR2HS $T=695640 628440 1 0 $X=695640 $Y=623020
X2279 2662 2651 2739 2 1 XNR2HS $T=699980 598200 0 0 $X=699980 $Y=597820
X2280 2740 2692 2726 2 1 XNR2HS $T=705560 678840 0 180 $X=699980 $Y=673420
X2281 2724 2729 2740 2 1 XNR2HS $T=699980 688920 1 0 $X=699980 $Y=683500
X2282 2631 2662 2749 2 1 XNR2HS $T=701220 628440 0 0 $X=701220 $Y=628060
X2283 2721 2753 2738 2 1 XNR2HS $T=707420 668760 1 180 $X=701840 $Y=668380
X2284 2747 2751 2754 2 1 XNR2HS $T=703700 567960 0 0 $X=703700 $Y=567580
X2285 2710 373 2773 2 1 XNR2HS $T=704940 688920 0 0 $X=704940 $Y=688540
X2286 2733 371 2767 2 1 XNR2HS $T=704940 709080 0 0 $X=704940 $Y=708700
X2287 2673 2765 2760 2 1 XNR2HS $T=711760 588120 1 180 $X=706180 $Y=587740
X2288 2631 2765 2784 2 1 XNR2HS $T=707420 618360 0 0 $X=707420 $Y=617980
X2289 2814 2810 2783 2 1 XNR2HS $T=715480 557880 1 180 $X=709900 $Y=557500
X2290 2782 2702 2790 2 1 XNR2HS $T=709900 567960 1 0 $X=709900 $Y=562540
X2291 369 374 2813 2 1 XNR2HS $T=710520 719160 1 0 $X=710520 $Y=713740
X2292 2790 2783 2818 2 1 XNR2HS $T=711140 557880 1 0 $X=711140 $Y=552460
X2293 2710 376 2793 2 1 XNR2HS $T=711140 688920 0 0 $X=711140 $Y=688540
X2294 2807 2738 2828 2 1 XNR2HS $T=712380 668760 1 0 $X=712380 $Y=663340
X2295 2845 2816 2819 2 1 XNR2HS $T=719200 648600 1 180 $X=713620 $Y=648220
X2296 2645 2631 2848 2 1 XNR2HS $T=714860 628440 0 0 $X=714860 $Y=628060
X2297 2823 2828 2833 2 1 XNR2HS $T=721060 658680 1 180 $X=715480 $Y=658300
X2298 2830 382 2851 2 1 XNR2HS $T=716100 699000 0 0 $X=716100 $Y=698620
X2299 2799 2630 2859 2 1 XNR2HS $T=716720 638520 1 0 $X=716720 $Y=633100
X2300 2830 389 2831 2 1 XNR2HS $T=722300 699000 0 180 $X=716720 $Y=693580
X2301 2720 2857 2869 2 1 XNR2HS $T=717960 598200 1 0 $X=717960 $Y=592780
X2302 2832 2875 2845 2 1 XNR2HS $T=724160 638520 1 180 $X=718580 $Y=638140
X2303 2849 2869 2894 2 1 XNR2HS $T=721060 588120 1 0 $X=721060 $Y=582700
X2304 2830 392 2880 2 1 XNR2HS $T=727880 699000 0 180 $X=722300 $Y=693580
X2305 2833 2888 2919 2 1 XNR2HS $T=723540 658680 1 0 $X=723540 $Y=653260
X2306 2808 2942 2924 2 1 XNR2HS $T=732840 567960 0 180 $X=727260 $Y=562540
X2307 2799 2685 2947 2 1 XNR2HS $T=727880 638520 1 0 $X=727880 $Y=633100
X2308 2630 2837 2955 2 1 XNR2HS $T=728500 618360 0 0 $X=728500 $Y=617980
X2309 2830 402 2914 2 1 XNR2HS $T=734080 699000 0 180 $X=728500 $Y=693580
X2310 2894 2936 403 2 1 XNR2HS $T=729740 557880 1 0 $X=729740 $Y=552460
X2311 2928 2944 2961 2 1 XNR2HS $T=729740 658680 1 0 $X=729740 $Y=653260
X2312 2986 2719 2843 2 1 XNR2HS $T=737800 578040 1 180 $X=732220 $Y=577660
X2313 2966 2934 2969 2 1 XNR2HS $T=739040 557880 1 180 $X=733460 $Y=557500
X2314 2967 2903 2990 2 1 XNR2HS $T=733460 668760 0 0 $X=733460 $Y=668380
X2315 2799 2719 2983 2 1 XNR2HS $T=734080 638520 1 0 $X=734080 $Y=633100
X2316 2981 2969 2998 2 1 XNR2HS $T=735320 557880 1 0 $X=735320 $Y=552460
X2317 3008 2762 2972 2 1 XNR2HS $T=740900 638520 1 180 $X=735320 $Y=638140
X2318 2973 396 2967 2 1 XNR2HS $T=735320 678840 1 0 $X=735320 $Y=673420
X2319 2987 2719 2976 2 1 XNR2HS $T=735940 598200 0 0 $X=735940 $Y=597820
X2320 2956 2961 3020 2 1 XNR2HS $T=737800 648600 0 0 $X=737800 $Y=648220
X2321 2792 2986 2984 2 1 XNR2HS $T=738420 578040 0 0 $X=738420 $Y=577660
X2322 3031 384 3010 2 1 XNR2HS $T=744620 668760 1 180 $X=739040 $Y=668380
X2323 2844 3009 3003 2 1 XNR2HS $T=739660 567960 1 0 $X=739660 $Y=562540
X2324 3008 2624 2989 2 1 XNR2HS $T=741520 618360 1 0 $X=741520 $Y=612940
X2325 2987 2715 3040 2 1 XNR2HS $T=749580 598200 1 180 $X=744000 $Y=597820
X2326 2988 3020 3060 2 1 XNR2HS $T=744000 648600 0 0 $X=744000 $Y=648220
X2327 402 2921 3043 2 1 XNR2HS $T=744000 699000 1 0 $X=744000 $Y=693580
X2328 3010 3047 3065 2 1 XNR2HS $T=744620 668760 0 0 $X=744620 $Y=668380
X2329 2649 3008 3038 2 1 XNR2HS $T=745240 638520 0 0 $X=745240 $Y=638140
X2330 3050 2935 3073 2 1 XNR2HS $T=745860 557880 1 0 $X=745860 $Y=552460
X2331 2715 3008 3056 2 1 XNR2HS $T=747100 648600 1 0 $X=747100 $Y=643180
X2332 3034 2978 3089 2 1 XNR2HS $T=749580 567960 0 0 $X=749580 $Y=567580
X2333 2986 2636 3096 2 1 XNR2HS $T=749580 578040 0 0 $X=749580 $Y=577660
X2334 3074 2636 3097 2 1 XNR2HS $T=749580 598200 0 0 $X=749580 $Y=597820
X2335 3048 2913 3098 2 1 XNR2HS $T=749580 658680 0 0 $X=749580 $Y=658300
X2336 415 3080 3099 2 1 XNR2HS $T=749580 678840 1 0 $X=749580 $Y=673420
X2337 3074 2624 3083 2 1 XNR2HS $T=755780 608280 0 180 $X=750200 $Y=602860
X2338 3077 3089 420 2 1 XNR2HS $T=750820 557880 0 0 $X=750820 $Y=557500
X2339 3068 389 3106 2 1 XNR2HS $T=750820 709080 1 0 $X=750820 $Y=703660
X2340 3073 3037 421 2 1 XNR2HS $T=751440 557880 1 0 $X=751440 $Y=552460
X2341 3074 2649 3115 2 1 XNR2HS $T=752680 618360 0 0 $X=752680 $Y=617980
X2342 3064 3079 3116 2 1 XNR2HS $T=752680 648600 1 0 $X=752680 $Y=643180
X2343 2624 2986 3129 2 1 XNR2HS $T=755160 578040 0 0 $X=755160 $Y=577660
X2344 2904 3099 3131 2 1 XNR2HS $T=755160 678840 1 0 $X=755160 $Y=673420
X2345 3139 3108 3119 2 1 XNR2HS $T=761980 547800 1 180 $X=756400 $Y=547420
X2346 3110 3098 3140 2 1 XNR2HS $T=756400 658680 0 0 $X=756400 $Y=658300
X2347 3068 392 3141 2 1 XNR2HS $T=756400 709080 1 0 $X=756400 $Y=703660
X2348 3036 3122 3145 2 1 XNR2HS $T=757020 668760 0 0 $X=757020 $Y=668380
X2349 3148 3144 3128 2 1 XNR2HS $T=763220 557880 0 180 $X=757640 $Y=552460
X2350 3086 3116 3149 2 1 XNR2HS $T=758880 648600 1 0 $X=758880 $Y=643180
X2351 3005 2762 3170 2 1 XNR2HS $T=761980 598200 0 0 $X=761980 $Y=597820
X2352 2975 3133 3176 2 1 XNR2HS $T=763220 578040 1 0 $X=763220 $Y=572620
X2353 3055 3138 3182 2 1 XNR2HS $T=763840 678840 1 0 $X=763840 $Y=673420
X2354 3005 2649 3193 2 1 XNR2HS $T=765080 588120 0 0 $X=765080 $Y=587740
X2355 3176 3184 3199 2 1 XNR2HS $T=766320 557880 1 0 $X=766320 $Y=552460
X2356 3164 3076 3204 2 1 XNR2HS $T=766940 628440 0 0 $X=766940 $Y=628060
X2357 3068 391 3206 2 1 XNR2HS $T=766940 719160 1 0 $X=766940 $Y=713740
X2358 3153 3145 3218 2 1 XNR2HS $T=768180 668760 0 0 $X=768180 $Y=668380
X2359 2839 3194 3227 2 1 XNR2HS $T=769420 688920 1 0 $X=769420 $Y=683500
X2360 3211 3199 3233 2 1 XNR2HS $T=770660 547800 0 0 $X=770660 $Y=547420
X2361 3239 3207 3221 2 1 XNR2HS $T=776860 557880 1 180 $X=771280 $Y=557500
X2362 2943 2785 3241 2 1 XNR2HS $T=771900 618360 0 0 $X=771900 $Y=617980
X2363 2802 3183 3243 2 1 XNR2HS $T=772520 699000 0 0 $X=772520 $Y=698620
X2364 3179 3085 3246 2 1 XNR2HS $T=773140 628440 0 0 $X=773140 $Y=628060
X2365 3209 3182 3256 2 1 XNR2HS $T=774380 678840 1 0 $X=774380 $Y=673420
X2366 3169 3067 3261 2 1 XNR2HS $T=775000 598200 1 0 $X=775000 $Y=592780
X2367 3246 3231 3266 2 1 XNR2HS $T=775620 638520 1 0 $X=775620 $Y=633100
X2368 3241 3156 3276 2 1 XNR2HS $T=777480 618360 0 0 $X=777480 $Y=617980
X2369 3088 3215 3277 2 1 XNR2HS $T=777480 688920 0 0 $X=777480 $Y=688540
X2370 3221 3196 3286 2 1 XNR2HS $T=778720 557880 1 0 $X=778720 $Y=552460
X2371 3304 3297 3280 2 1 XNR2HS $T=786160 557880 1 180 $X=780580 $Y=557500
X2372 3114 3084 3298 2 1 XNR2HS $T=780580 598200 0 0 $X=780580 $Y=597820
X2373 3107 3270 3305 2 1 XNR2HS $T=781820 588120 0 0 $X=781820 $Y=587740
X2374 3251 3147 3306 2 1 XNR2HS $T=781820 628440 1 0 $X=781820 $Y=623020
X2375 3227 3284 3308 2 1 XNR2HS $T=781820 688920 1 0 $X=781820 $Y=683500
X2376 3290 3261 3297 2 1 XNR2HS $T=788640 567960 0 180 $X=783060 $Y=562540
X2377 3219 3277 3291 2 1 XNR2HS $T=783060 688920 0 0 $X=783060 $Y=688540
X2378 3032 3272 3317 2 1 XNR2HS $T=783680 709080 1 0 $X=783680 $Y=703660
X2379 3103 3263 3324 2 1 XNR2HS $T=784920 699000 0 0 $X=784920 $Y=698620
X2380 2840 3174 3325 2 1 XNR2HS $T=784920 709080 0 0 $X=784920 $Y=708700
X2381 3001 3259 3335 2 1 XNR2HS $T=786780 719160 1 0 $X=786780 $Y=713740
X2382 3224 3305 3319 2 1 XNR2HS $T=787400 588120 0 0 $X=787400 $Y=587740
X2383 3291 3308 3338 2 1 XNR2HS $T=787400 688920 1 0 $X=787400 $Y=683500
X2384 3210 3324 3342 2 1 XNR2HS $T=788020 699000 1 0 $X=788020 $Y=693580
X2385 3242 3292 3349 2 1 XNR2HS $T=788640 688920 0 0 $X=788640 $Y=688540
X2386 3317 3258 3352 2 1 XNR2HS $T=789260 709080 1 0 $X=789260 $Y=703660
X2387 3298 3312 3366 2 1 XNR2HS $T=791120 578040 0 0 $X=791120 $Y=577660
X2388 3341 3307 3374 2 1 XNR2HS $T=792360 628440 0 0 $X=792360 $Y=628060
X2389 3243 3369 3392 2 1 XNR2HS $T=794840 709080 1 0 $X=794840 $Y=703660
X2390 3352 3392 3413 2 1 XNR2HS $T=798560 699000 0 0 $X=798560 $Y=698620
X2391 441 3335 3414 2 1 XNR2HS $T=798560 719160 1 0 $X=798560 $Y=713740
X2392 3349 3342 3417 2 1 XNR2HS $T=799180 688920 0 0 $X=799180 $Y=688540
X2393 3385 3410 448 2 1 XNR2HS $T=802900 547800 0 0 $X=802900 $Y=547420
X2394 3519 3356 3536 2 1 XNR2HS $T=820260 678840 0 0 $X=820260 $Y=678460
X2395 461 463 3532 2 1 XNR2HS $T=821500 709080 0 0 $X=821500 $Y=708700
X2396 3452 3549 3559 2 1 XNR2HS $T=826460 678840 0 0 $X=826460 $Y=678460
X2397 3533 3554 3574 2 1 XNR2HS $T=829560 709080 1 0 $X=829560 $Y=703660
X2398 3557 3544 3577 2 1 XNR2HS $T=830180 699000 0 0 $X=830180 $Y=698620
X2399 3421 3572 3590 2 1 XNR2HS $T=832040 668760 1 0 $X=832040 $Y=663340
X2400 3586 3591 3607 2 1 XNR2HS $T=835760 678840 1 0 $X=835760 $Y=673420
X2401 3598 3579 3648 2 1 XNR2HS $T=842580 618360 1 0 $X=842580 $Y=612940
X2402 3628 3584 3658 2 1 XNR2HS $T=843820 618360 0 0 $X=843820 $Y=617980
X2403 3728 3724 3712 2 1 XNR2HS $T=867380 638520 1 180 $X=861800 $Y=638140
X2404 3741 3733 3717 2 1 XNR2HS $T=869240 648600 0 180 $X=863660 $Y=643180
X2405 3790 3787 3721 2 1 XNR2HS $T=877920 638520 0 180 $X=872340 $Y=633100
X2406 3829 3807 3808 2 1 XNR2HS $T=884120 628440 1 180 $X=878540 $Y=628060
X2407 525 3834 3788 2 1 XNR2HS $T=885360 719160 0 180 $X=879780 $Y=713740
X2408 530 529 3834 2 1 XNR2HS $T=888460 709080 1 180 $X=882880 $Y=708700
X2409 3869 3853 3842 2 1 XNR2HS $T=890940 628440 1 180 $X=885360 $Y=628060
X2410 3873 3866 3848 2 1 XNR2HS $T=891560 688920 0 180 $X=885980 $Y=683500
X2411 3856 3827 3871 2 1 XNR2HS $T=886600 547800 1 0 $X=886600 $Y=542380
X2412 3747 533 3895 2 1 XNR2HS $T=890320 547800 0 0 $X=890320 $Y=547420
X2413 3912 3862 3886 2 1 XNR2HS $T=897140 678840 1 180 $X=891560 $Y=678460
X2414 3772 3879 3907 2 1 XNR2HS $T=892180 557880 1 0 $X=892180 $Y=552460
X2415 3924 3918 3851 2 1 XNR2HS $T=899000 628440 1 180 $X=893420 $Y=628060
X2416 3925 3920 3893 2 1 XNR2HS $T=899000 709080 0 180 $X=893420 $Y=703660
X2417 3904 3917 3936 2 1 XNR2HS $T=895900 598200 1 0 $X=895900 $Y=592780
X2418 3890 3926 3955 2 1 XNR2HS $T=898380 557880 1 0 $X=898380 $Y=552460
X2419 549 3963 3920 2 1 XNR2HS $T=905200 709080 0 180 $X=899620 $Y=703660
X2420 3948 3931 3940 2 1 XNR2HS $T=900240 628440 0 0 $X=900240 $Y=628060
X2421 554 3988 3925 2 1 XNR2HS $T=909540 719160 0 180 $X=903960 $Y=713740
X2422 3993 3987 4008 2 1 XNR2HS $T=907680 638520 1 0 $X=907680 $Y=633100
X2423 563 559 3988 2 1 XNR2HS $T=915740 719160 0 180 $X=910160 $Y=713740
X2424 4050 4031 4024 2 1 XNR2HS $T=918840 699000 1 180 $X=913260 $Y=698620
X2425 4051 566 4031 2 1 XNR2HS $T=918840 709080 0 180 $X=913260 $Y=703660
X2426 4074 4069 4054 2 1 XNR2HS $T=922560 638520 0 180 $X=916980 $Y=633100
X2427 571 570 4050 2 1 XNR2HS $T=923800 719160 0 180 $X=918220 $Y=713740
X2428 4065 4067 4089 2 1 XNR2HS $T=919460 678840 1 0 $X=919460 $Y=673420
X2429 4104 4098 4073 2 1 XNR2HS $T=925660 628440 0 180 $X=920080 $Y=623020
X2430 4085 4093 4106 2 1 XNR2HS $T=921940 699000 1 0 $X=921940 $Y=693580
X2431 575 574 4051 2 1 XNR2HS $T=930000 709080 1 180 $X=924420 $Y=708700
X2432 4144 4122 4121 2 1 XNR2HS $T=932480 618360 1 180 $X=926900 $Y=617980
X2433 576 577 4093 2 1 XNR2HS $T=933100 699000 0 180 $X=927520 $Y=693580
X2434 578 4146 4085 2 1 XNR2HS $T=933720 709080 0 180 $X=928140 $Y=703660
X2435 582 4143 4146 2 1 XNR2HS $T=937440 719160 0 180 $X=931860 $Y=713740
X2436 4169 4163 4181 2 1 XNR2HS $T=938060 628440 1 0 $X=938060 $Y=623020
X2437 586 590 4186 2 1 XNR2HS $T=938680 719160 1 0 $X=938680 $Y=713740
X2438 4176 4129 4189 2 1 XNR2HS $T=939300 678840 0 0 $X=939300 $Y=678460
X2439 594 595 4217 2 1 XNR2HS $T=947360 719160 1 0 $X=947360 $Y=713740
X2440 4256 4254 4265 2 1 XNR2HS $T=961000 678840 1 0 $X=961000 $Y=673420
X2441 1057 841 1084 1 2 XOR2H $T=337900 588120 0 0 $X=337900 $Y=587740
X2442 92 86 81 1 2 XOR2H $T=409820 719160 0 180 $X=401140 $Y=713740
X2443 3195 3354 3389 1 2 XOR2H $T=791740 638520 0 0 $X=791740 $Y=638140
X2444 3514 3509 454 1 2 XOR2H $T=819640 608280 0 180 $X=810960 $Y=602860
X2445 695 2 721 697 1 NR2 $T=274660 648600 1 0 $X=274660 $Y=643180
X2446 767 2 781 739 1 NR2 $T=285820 578040 1 0 $X=285820 $Y=572620
X2447 780 2 759 774 1 NR2 $T=288920 668760 1 180 $X=287060 $Y=668380
X2448 767 2 769 785 1 NR2 $T=289540 567960 0 0 $X=289540 $Y=567580
X2449 785 2 804 781 1 NR2 $T=291400 578040 0 180 $X=289540 $Y=572620
X2450 828 2 835 837 1 NR2 $T=297600 668760 0 0 $X=297600 $Y=668380
X2451 865 2 900 889 1 NR2 $T=308140 547800 0 0 $X=308140 $Y=547420
X2452 894 2 882 901 1 NR2 $T=308760 608280 0 0 $X=308760 $Y=607900
X2453 884 2 923 913 1 NR2 $T=314340 557880 1 0 $X=314340 $Y=552460
X2454 900 2 22 923 1 NR2 $T=316820 547800 0 0 $X=316820 $Y=547420
X2455 909 2 954 940 1 NR2 $T=319300 567960 1 0 $X=319300 $Y=562540
X2456 955 2 968 949 1 NR2 $T=321160 628440 0 180 $X=319300 $Y=623020
X2457 816 2 31 990 1 NR2 $T=329840 547800 1 0 $X=329840 $Y=542380
X2458 973 2 1044 1032 1 NR2 $T=335420 557880 0 0 $X=335420 $Y=557500
X2459 1000 2 1029 1042 1 NR2 $T=339140 608280 1 0 $X=339140 $Y=602860
X2460 1041 2 1085 943 1 NR2 $T=344100 567960 1 0 $X=344100 $Y=562540
X2461 1074 2 1126 1008 1 NR2 $T=349680 557880 0 0 $X=349680 $Y=557500
X2462 1143 2 1148 1128 1 NR2 $T=354640 578040 0 180 $X=352780 $Y=572620
X2463 954 2 1152 1085 1 NR2 $T=353400 567960 0 0 $X=353400 $Y=567580
X2464 1173 2 1090 1179 1 NR2 $T=359600 628440 0 0 $X=359600 $Y=628060
X2465 1134 2 53 1113 1 NR2 $T=360220 547800 1 0 $X=360220 $Y=542380
X2466 1044 2 1172 1126 1 NR2 $T=360220 557880 0 0 $X=360220 $Y=557500
X2467 918 2 1188 1175 1 NR2 $T=362700 618360 0 180 $X=360840 $Y=612940
X2468 1171 2 1135 1220 1 NR2 $T=362700 557880 1 0 $X=362700 $Y=552460
X2469 1195 2 1137 1200 1 NR2 $T=362700 608280 0 0 $X=362700 $Y=607900
X2470 1173 2 874 1201 1 NR2 $T=362700 628440 0 0 $X=362700 $Y=628060
X2471 1085 2 1212 1208 1 NR2 $T=363940 567960 0 0 $X=363940 $Y=567580
X2472 1222 2 1204 1154 1 NR2 $T=366420 699000 0 180 $X=364560 $Y=693580
X2473 1228 2 919 1173 1 NR2 $T=367660 638520 0 180 $X=365800 $Y=633100
X2474 1218 2 58 1170 1 NR2 $T=367660 547800 1 0 $X=367660 $Y=542380
X2475 1230 2 1169 1243 1 NR2 $T=368900 608280 1 0 $X=368900 $Y=602860
X2476 53 2 1250 58 1 NR2 $T=369520 547800 1 0 $X=369520 $Y=542380
X2477 1271 2 1265 1266 1 NR2 $T=375720 618360 0 180 $X=373860 $Y=612940
X2478 1234 2 827 1295 1 NR2 $T=376960 638520 0 0 $X=376960 $Y=638140
X2479 1240 2 1300 1252 1 NR2 $T=378820 648600 1 180 $X=376960 $Y=648220
X2480 1315 2 1301 1234 1 NR2 $T=381920 638520 1 180 $X=380060 $Y=638140
X2481 1313 2 1276 1236 1 NR2 $T=381920 628440 1 0 $X=381920 $Y=623020
X2482 1316 2 1319 1262 1 NR2 $T=385640 547800 1 180 $X=383780 $Y=547420
X2483 1319 2 64 1336 1 NR2 $T=385020 547800 1 0 $X=385020 $Y=542380
X2484 1332 2 1261 1321 1 NR2 $T=385640 628440 0 0 $X=385640 $Y=628060
X2485 1341 2 1359 71 1 NR2 $T=388740 709080 1 0 $X=388740 $Y=703660
X2486 1360 2 1336 1374 1 NR2 $T=391220 547800 0 0 $X=391220 $Y=547420
X2487 1365 2 1353 1236 1 NR2 $T=393080 618360 1 180 $X=391220 $Y=617980
X2488 1295 2 1372 1202 1 NR2 $T=394320 638520 0 180 $X=392460 $Y=633100
X2489 1362 2 1388 1323 1 NR2 $T=395560 588120 0 180 $X=393700 $Y=582700
X2490 1357 2 1363 1368 1 NR2 $T=397420 608280 0 0 $X=397420 $Y=607900
X2491 1391 2 1329 786 1 NR2 $T=399900 648600 0 0 $X=399900 $Y=648220
X2492 1410 2 1397 1420 1 NR2 $T=401140 608280 0 0 $X=401140 $Y=607900
X2493 1228 2 1405 1436 1 NR2 $T=403000 648600 1 0 $X=403000 $Y=643180
X2494 1315 2 1435 786 1 NR2 $T=407340 638520 0 180 $X=405480 $Y=633100
X2495 1439 2 1384 1447 1 NR2 $T=407340 638520 1 0 $X=407340 $Y=633100
X2496 1438 2 1427 1442 1 NR2 $T=409820 688920 0 0 $X=409820 $Y=688540
X2497 1472 2 1448 1453 1 NR2 $T=413540 648600 1 0 $X=413540 $Y=643180
X2498 1295 2 1506 1443 1 NR2 $T=420360 618360 0 180 $X=418500 $Y=612940
X2499 1382 2 1510 1315 1 NR2 $T=418500 638520 0 0 $X=418500 $Y=638140
X2500 101 2 1479 1509 1 NR2 $T=419740 709080 1 0 $X=419740 $Y=703660
X2501 1505 2 1522 1441 1 NR2 $T=422840 678840 0 180 $X=420980 $Y=673420
X2502 1500 2 1441 1486 1 NR2 $T=422840 678840 0 0 $X=422840 $Y=678460
X2503 1523 2 1494 108 1 NR2 $T=424080 709080 1 0 $X=424080 $Y=703660
X2504 105 2 1531 1516 1 NR2 $T=429660 699000 0 0 $X=429660 $Y=698620
X2505 1564 2 1571 1548 1 NR2 $T=432760 608280 1 180 $X=430900 $Y=607900
X2506 1499 2 1556 1240 1 NR2 $T=433380 628440 1 180 $X=431520 $Y=628060
X2507 1515 2 1570 1475 1 NR2 $T=432140 598200 1 0 $X=432140 $Y=592780
X2508 1559 2 1558 1552 1 NR2 $T=432140 688920 1 0 $X=432140 $Y=683500
X2509 1574 2 1572 1560 1 NR2 $T=435860 618360 0 180 $X=434000 $Y=612940
X2510 1499 2 1578 1267 1 NR2 $T=437100 628440 1 180 $X=435240 $Y=628060
X2511 1435 2 1605 1433 1 NR2 $T=436480 638520 1 0 $X=436480 $Y=633100
X2512 1584 2 1503 118 1 NR2 $T=436480 709080 1 0 $X=436480 $Y=703660
X2513 1593 2 1595 1558 1 NR2 $T=438960 668760 1 180 $X=437100 $Y=668380
X2514 1571 2 1612 1572 1 NR2 $T=439580 608280 1 0 $X=439580 $Y=602860
X2515 1626 2 1614 1611 1 NR2 $T=443300 688920 1 180 $X=441440 $Y=688540
X2516 1622 2 1620 1615 1 NR2 $T=445780 618360 1 180 $X=443920 $Y=617980
X2517 1556 2 1627 1625 1 NR2 $T=443920 628440 0 0 $X=443920 $Y=628060
X2518 1640 2 1655 1620 1 NR2 $T=449500 618360 0 0 $X=449500 $Y=617980
X2519 131 2 1651 1667 1 NR2 $T=453220 709080 0 0 $X=453220 $Y=708700
X2520 1656 2 1681 1662 1 NR2 $T=454460 638520 1 0 $X=454460 $Y=633100
X2521 1651 2 1671 1649 1 NR2 $T=454460 699000 1 0 $X=454460 $Y=693580
X2522 1671 2 1683 1659 1 NR2 $T=456940 688920 0 0 $X=456940 $Y=688540
X2523 115 2 1707 1394 1 NR2 $T=458800 719160 0 180 $X=456940 $Y=713740
X2524 1669 2 1686 1450 1 NR2 $T=458180 547800 0 0 $X=458180 $Y=547420
X2525 1666 2 1670 1703 1 NR2 $T=460040 709080 1 0 $X=460040 $Y=703660
X2526 1704 2 1700 1670 1 NR2 $T=462520 699000 1 180 $X=460660 $Y=698620
X2527 1707 2 1719 136 1 NR2 $T=463140 719160 1 0 $X=463140 $Y=713740
X2528 1701 2 1713 1695 1 NR2 $T=464380 578040 1 0 $X=464380 $Y=572620
X2529 1686 2 1730 1731 1 NR2 $T=466240 557880 1 0 $X=466240 $Y=552460
X2530 1708 2 1731 1706 1 NR2 $T=468100 557880 1 180 $X=466240 $Y=557500
X2531 142 2 1749 1729 1 NR2 $T=467480 618360 1 0 $X=467480 $Y=612940
X2532 1702 2 1743 1733 1 NR2 $T=468720 598200 1 0 $X=468720 $Y=592780
X2533 147 2 1716 1728 1 NR2 $T=470580 719160 0 180 $X=468720 $Y=713740
X2534 1712 2 1773 1735 1 NR2 $T=472440 578040 0 0 $X=472440 $Y=577660
X2535 1697 2 1777 1685 1 NR2 $T=472440 588120 0 0 $X=472440 $Y=587740
X2536 1734 2 1781 1760 1 NR2 $T=473680 608280 1 0 $X=473680 $Y=602860
X2537 1713 2 1772 1773 1 NR2 $T=474300 567960 0 0 $X=474300 $Y=567580
X2538 1777 2 1785 1743 1 NR2 $T=476160 588120 0 0 $X=476160 $Y=587740
X2539 1731 2 1795 1780 1 NR2 $T=479880 567960 0 180 $X=478020 $Y=562540
X2540 2639 2 2635 2628 1 NR2 $T=683240 618360 1 180 $X=681380 $Y=617980
X2541 2674 2 359 2666 1 NR2 $T=691920 557880 0 180 $X=690060 $Y=552460
X2542 2678 2 2669 2663 1 NR2 $T=692540 588120 0 180 $X=690680 $Y=582700
X2543 2669 2 2686 2681 1 NR2 $T=691920 578040 0 0 $X=691920 $Y=577660
X2544 2687 2 2689 2638 1 NR2 $T=695020 608280 0 180 $X=693160 $Y=602860
X2545 2688 2 2694 2699 1 NR2 $T=695640 578040 0 0 $X=695640 $Y=577660
X2546 2694 2 2670 2675 1 NR2 $T=696260 567960 1 0 $X=696260 $Y=562540
X2547 2682 2 2707 2687 1 NR2 $T=701220 628440 1 180 $X=699360 $Y=628060
X2548 2716 2 2732 2730 1 NR2 $T=699980 547800 0 0 $X=699980 $Y=547420
X2549 2734 2 363 2705 1 NR2 $T=703080 557880 1 180 $X=701220 $Y=557500
X2550 2735 2 368 2688 1 NR2 $T=703080 578040 0 180 $X=701220 $Y=572620
X2551 372 2 2708 2731 1 NR2 $T=704320 709080 0 180 $X=702460 $Y=703660
X2552 2746 2 2716 2771 1 NR2 $T=706180 547800 0 0 $X=706180 $Y=547420
X2553 2755 2 2785 2682 1 NR2 $T=708660 638520 1 0 $X=708660 $Y=633100
X2554 2682 2 2795 2778 1 NR2 $T=711140 638520 0 0 $X=711140 $Y=638140
X2555 2797 2 2711 2680 1 NR2 $T=713620 578040 0 180 $X=711760 $Y=572620
X2556 2765 2 2797 2825 1 NR2 $T=712380 588120 0 0 $X=712380 $Y=587740
X2557 2826 2 2822 2745 1 NR2 $T=715480 628440 0 180 $X=713620 $Y=623020
X2558 2604 2 2798 2829 1 NR2 $T=714240 618360 1 0 $X=714240 $Y=612940
X2559 2736 2 2853 2825 1 NR2 $T=716100 578040 0 0 $X=716100 $Y=577660
X2560 2765 2 2841 2826 1 NR2 $T=717340 618360 0 0 $X=717340 $Y=617980
X2561 2851 2 2864 2838 1 NR2 $T=719200 678840 1 180 $X=717340 $Y=678460
X2562 2826 2 2878 2805 1 NR2 $T=720440 618360 1 0 $X=720440 $Y=612940
X2563 2867 2 2882 2864 1 NR2 $T=721060 678840 0 0 $X=721060 $Y=678460
X2564 2805 2 2861 2872 1 NR2 $T=723540 618360 1 0 $X=723540 $Y=612940
X2565 2749 2 2895 2884 1 NR2 $T=724160 628440 1 0 $X=724160 $Y=623020
X2566 390 2 2911 2915 1 NR2 $T=725400 719160 1 0 $X=725400 $Y=713740
X2567 2709 2 2932 2887 1 NR2 $T=727880 628440 1 180 $X=726020 $Y=628060
X2568 2872 2 2931 2709 1 NR2 $T=729120 628440 0 180 $X=727260 $Y=623020
X2569 367 2 397 2911 1 NR2 $T=727880 719160 1 0 $X=727880 $Y=713740
X2570 2931 2 2935 2895 1 NR2 $T=731600 628440 0 180 $X=729740 $Y=623020
X2571 2942 2 2981 2982 1 NR2 $T=734700 567960 1 0 $X=734700 $Y=562540
X2572 2912 2 2964 2848 1 NR2 $T=736560 628440 1 180 $X=734700 $Y=628060
X2573 2949 2 2948 2921 1 NR2 $T=735320 699000 1 0 $X=735320 $Y=693580
X2574 2956 2 2997 2961 1 NR2 $T=735940 658680 1 0 $X=735940 $Y=653260
X2575 2935 2 3054 3063 1 NR2 $T=745240 557880 0 0 $X=745240 $Y=557500
X2576 3009 2 3077 3051 1 NR2 $T=747720 567960 1 0 $X=747720 $Y=562540
X2577 3073 2 3082 3037 1 NR2 $T=750200 547800 0 0 $X=750200 $Y=547420
X2578 3064 2 3104 3086 1 NR2 $T=757640 648600 0 0 $X=757640 $Y=648220
X2579 3133 2 3146 3117 1 NR2 $T=761980 578040 0 180 $X=760120 $Y=572620
X2580 3142 2 3153 2882 1 NR2 $T=763220 678840 0 180 $X=761360 $Y=673420
X2581 2788 2 3158 2898 1 NR2 $T=763220 658680 0 0 $X=763220 $Y=658300
X2582 3139 2 3168 3108 1 NR2 $T=765700 557880 0 180 $X=763840 $Y=552460
X2583 3166 2 3178 3156 1 NR2 $T=767560 618360 1 180 $X=765700 $Y=617980
X2584 3155 2 3279 3149 1 NR2 $T=771900 648600 1 180 $X=770040 $Y=648220
X2585 3183 2 3210 3188 1 NR2 $T=772520 699000 1 180 $X=770660 $Y=698620
X2586 3194 2 3209 3205 1 NR2 $T=771280 678840 0 0 $X=771280 $Y=678460
X2587 3157 2 3269 3016 1 NR2 $T=779340 588120 0 0 $X=779340 $Y=587740
X2588 3227 2 3288 3284 1 NR2 $T=780580 678840 1 0 $X=780580 $Y=673420
X2589 3174 2 3272 3285 1 NR2 $T=780580 709080 0 0 $X=780580 $Y=708700
X2590 3114 2 3299 3271 1 NR2 $T=781200 608280 0 0 $X=781200 $Y=607900
X2591 3261 2 3294 3290 1 NR2 $T=781820 567960 0 0 $X=781820 $Y=567580
X2592 3150 2 3300 3252 1 NR2 $T=785540 648600 0 180 $X=783680 $Y=643180
X2593 3280 2 3339 3283 1 NR2 $T=791120 557880 0 0 $X=791120 $Y=557500
X2594 3243 2 3368 3369 1 NR2 $T=795460 699000 0 0 $X=795460 $Y=698620
X2595 2985 2 3418 3333 1 NR2 $T=801040 638520 1 0 $X=801040 $Y=633100
X2596 3409 2 3442 3338 1 NR2 $T=802900 688920 1 0 $X=802900 $Y=683500
X2597 3430 2 3444 3408 1 NR2 $T=804140 678840 0 0 $X=804140 $Y=678460
X2598 3413 2 3485 3428 1 NR2 $T=811580 699000 0 180 $X=809720 $Y=693580
X2599 3525 2 3533 3466 1 NR2 $T=822740 709080 0 180 $X=820880 $Y=703660
X2600 466 2 3542 2223 1 NR2 $T=823980 618360 0 0 $X=823980 $Y=617980
X2601 3583 2 3589 3529 1 NR2 $T=833900 588120 1 180 $X=832040 $Y=587740
X2602 3566 2 3609 3552 1 NR2 $T=837620 608280 0 180 $X=835760 $Y=602860
X2603 471 2 3597 473 1 NR2 $T=836380 709080 0 0 $X=836380 $Y=708700
X2604 476 2 3596 3604 1 NR2 $T=839480 709080 1 0 $X=839480 $Y=703660
X2605 3596 2 3622 3597 1 NR2 $T=840100 688920 0 0 $X=840100 $Y=688540
X2606 3594 2 3651 3565 1 NR2 $T=843200 567960 0 0 $X=843200 $Y=567580
X2607 3619 2 3633 3640 1 NR2 $T=843200 578040 0 0 $X=843200 $Y=577660
X2608 485 2 3626 486 1 NR2 $T=846920 547800 1 180 $X=845060 $Y=547420
X2609 3636 2 3659 3539 1 NR2 $T=845680 598200 1 0 $X=845680 $Y=592780
X2610 3599 2 3650 3623 1 NR2 $T=845680 709080 1 0 $X=845680 $Y=703660
X2611 480 2 3667 488 1 NR2 $T=846300 547800 1 0 $X=846300 $Y=542380
X2612 3651 2 3653 3633 1 NR2 $T=846300 567960 0 0 $X=846300 $Y=567580
X2613 3650 2 3654 3632 1 NR2 $T=848160 678840 0 180 $X=846300 $Y=673420
X2614 3635 2 3617 3650 1 NR2 $T=848160 699000 0 180 $X=846300 $Y=693580
X2615 3655 2 3635 3671 1 NR2 $T=846920 699000 0 0 $X=846920 $Y=698620
X2616 3589 2 3675 3659 1 NR2 $T=848160 588120 0 0 $X=848160 $Y=587740
X2617 3667 2 3660 3626 1 NR2 $T=853740 547800 1 180 $X=851880 $Y=547420
X2618 3687 2 3692 3664 1 NR2 $T=853740 557880 0 180 $X=851880 $Y=552460
X2619 3626 2 3687 3686 1 NR2 $T=852500 557880 0 0 $X=852500 $Y=557500
X2620 3715 2 502 3723 1 NR2 $T=863040 719160 1 0 $X=863040 $Y=713740
X2621 3738 2 506 504 1 NR2 $T=865520 547800 0 180 $X=863660 $Y=542380
X2622 3710 2 3730 3739 1 NR2 $T=866140 557880 0 0 $X=866140 $Y=557500
X2623 3708 2 3731 3729 1 NR2 $T=866760 658680 0 0 $X=866760 $Y=658300
X2624 3762 2 3746 3731 1 NR2 $T=871720 648600 1 180 $X=869860 $Y=648220
X2625 3767 2 3735 3749 1 NR2 $T=872340 709080 0 180 $X=870480 $Y=703660
X2626 3774 2 3762 3763 1 NR2 $T=872960 668760 0 180 $X=871100 $Y=663340
X2627 3740 2 3751 3765 1 NR2 $T=873580 578040 0 0 $X=873580 $Y=577660
X2628 3751 2 3769 3784 1 NR2 $T=874200 557880 0 0 $X=874200 $Y=557500
X2629 3784 2 3795 3782 1 NR2 $T=877300 557880 0 180 $X=875440 $Y=552460
X2630 3730 2 3776 520 1 NR2 $T=876680 547800 1 0 $X=876680 $Y=542380
X2631 3720 2 3784 3779 1 NR2 $T=879160 567960 1 180 $X=877300 $Y=567580
X2632 3793 2 3796 3806 1 NR2 $T=877300 578040 0 0 $X=877300 $Y=577660
X2633 3800 2 3749 3820 1 NR2 $T=877920 709080 1 0 $X=877920 $Y=703660
X2634 3819 2 3811 3817 1 NR2 $T=882260 658680 1 180 $X=880400 $Y=658300
X2635 3791 2 3832 3816 1 NR2 $T=881020 588120 1 0 $X=881020 $Y=582700
X2636 3799 2 3817 3814 1 NR2 $T=881020 668760 1 0 $X=881020 $Y=663340
X2637 3804 2 3836 3821 1 NR2 $T=882260 567960 0 0 $X=882260 $Y=567580
X2638 3832 2 3846 3796 1 NR2 $T=884740 578040 1 180 $X=882880 $Y=577660
X2639 3843 2 3849 3833 1 NR2 $T=885360 648600 0 180 $X=883500 $Y=643180
X2640 3839 2 3819 3850 1 NR2 $T=884120 658680 0 0 $X=884120 $Y=658300
X2641 528 2 3877 3835 1 NR2 $T=889700 567960 1 0 $X=889700 $Y=562540
X2642 3865 2 3884 3872 1 NR2 $T=891560 658680 0 0 $X=891560 $Y=658300
X2643 3910 2 3885 3884 1 NR2 $T=894040 658680 0 180 $X=892180 $Y=653260
X2644 3905 2 3898 3893 1 NR2 $T=895280 699000 0 180 $X=893420 $Y=693580
X2645 3836 2 3906 3877 1 NR2 $T=894660 567960 0 0 $X=894660 $Y=567580
X2646 3934 2 3910 3937 1 NR2 $T=898380 658680 0 0 $X=898380 $Y=658300
X2647 3927 2 3873 3945 1 NR2 $T=898380 688920 1 0 $X=898380 $Y=683500
X2648 3952 2 3891 3939 1 NR2 $T=902100 638520 1 180 $X=900240 $Y=638140
X2649 3953 2 3952 3968 1 NR2 $T=901480 658680 1 0 $X=901480 $Y=653260
X2650 3975 2 3932 3952 1 NR2 $T=903960 648600 1 180 $X=902100 $Y=648220
X2651 3972 2 3971 3956 1 NR2 $T=905820 578040 0 180 $X=903960 $Y=572620
X2652 3977 2 551 3956 1 NR2 $T=907060 567960 0 180 $X=905200 $Y=562540
X2653 3923 2 3972 4017 1 NR2 $T=911400 578040 1 0 $X=911400 $Y=572620
X2654 4011 2 3975 4000 1 NR2 $T=911400 658680 1 0 $X=911400 $Y=653260
X2655 4043 2 4042 4024 1 NR2 $T=916360 699000 1 0 $X=916360 $Y=693580
X2656 4068 2 4040 3901 1 NR2 $T=919460 557880 1 180 $X=917600 $Y=557500
X2657 4061 2 4046 4075 1 NR2 $T=919460 567960 1 0 $X=919460 $Y=562540
X2658 4064 2 4009 4081 1 NR2 $T=920080 638520 0 0 $X=920080 $Y=638140
X2659 3823 2 4076 4082 1 NR2 $T=921320 588120 0 0 $X=921320 $Y=587740
X2660 4084 2 4064 4037 1 NR2 $T=923180 648600 1 180 $X=921320 $Y=648220
X2661 4130 2 4113 4046 1 NR2 $T=928140 557880 0 180 $X=926280 $Y=552460
X2662 4087 2 4130 573 1 NR2 $T=926900 547800 0 0 $X=926900 $Y=547420
X2663 4099 2 4127 4078 1 NR2 $T=927520 598200 1 0 $X=927520 $Y=592780
X2664 4107 2 4143 575 1 NR2 $T=930000 719160 0 180 $X=928140 $Y=713740
X2665 4128 2 4083 4110 1 NR2 $T=930620 648600 0 180 $X=928760 $Y=643180
X2666 4118 2 4135 4083 1 NR2 $T=931240 638520 0 180 $X=929380 $Y=633100
X2667 4127 2 4105 4076 1 NR2 $T=930000 588120 1 0 $X=930000 $Y=582700
X2668 4145 2 4118 4151 1 NR2 $T=931860 648600 1 0 $X=931860 $Y=643180
X2669 4046 2 4136 4155 1 NR2 $T=934340 567960 1 0 $X=934340 $Y=562540
X2670 4177 2 4159 4165 1 NR2 $T=939300 638520 1 180 $X=937440 $Y=638140
X2671 4166 2 4165 4175 1 NR2 $T=937440 648600 1 0 $X=937440 $Y=643180
X2672 4172 2 4190 4154 1 NR2 $T=940540 699000 0 0 $X=940540 $Y=698620
X2673 4199 2 4177 4191 1 NR2 $T=949220 638520 1 180 $X=947360 $Y=638140
X2674 4167 2 4225 4219 1 NR2 $T=950460 547800 0 0 $X=950460 $Y=547420
X2675 4243 2 601 4225 1 NR2 $T=956040 547800 0 180 $X=954180 $Y=542380
X2676 4224 2 4243 4229 1 NR2 $T=955420 557880 1 0 $X=955420 $Y=552460
X2677 4227 2 4237 4207 1 NR2 $T=957900 688920 0 180 $X=956040 $Y=683500
X2678 4260 2 608 4263 1 NR2 $T=961620 547800 1 0 $X=961620 $Y=542380
X2679 4262 2 4263 4270 1 NR2 $T=962240 547800 0 0 $X=962240 $Y=547420
X2680 4283 2 4260 4305 1 NR2 $T=969060 547800 1 0 $X=969060 $Y=542380
X2681 618 2 4350 4352 1 NR2 $T=988900 699000 1 0 $X=988900 $Y=693580
X2682 623 2 4342 618 1 NR2 $T=988900 709080 0 0 $X=988900 $Y=708700
X2683 693 2 714 1 696 NR2P $T=266600 628440 0 180 $X=262880 $Y=623020
X2684 710 2 698 1 724 NR2P $T=269700 588120 1 180 $X=265980 $Y=587740
X2685 716 2 737 1 698 NR2P $T=271560 598200 0 180 $X=267840 $Y=592780
X2686 735 2 724 1 739 NR2P $T=272800 588120 0 0 $X=272800 $Y=587740
X2687 768 2 739 1 777 NR2P $T=283960 588120 0 0 $X=283960 $Y=587740
X2688 707 2 767 1 776 NR2P $T=288300 578040 1 180 $X=284580 $Y=577660
X2689 707 2 768 1 794 NR2P $T=290780 588120 0 180 $X=287060 $Y=582700
X2690 798 2 777 1 807 NR2P $T=290160 588120 0 0 $X=290160 $Y=587740
X2691 859 2 846 1 840 NR2P $T=301320 608280 1 0 $X=301320 $Y=602860
X2692 899 2 886 1 772 NR2P $T=307520 598200 1 0 $X=307520 $Y=592780
X2693 994 2 995 1 907 NR2P $T=326120 678840 0 0 $X=326120 $Y=678460
X2694 1033 2 1028 1 966 NR2P $T=332940 588120 1 0 $X=332940 $Y=582700
X2695 1049 2 1055 1 896 NR2P $T=334800 668760 0 0 $X=334800 $Y=668380
X2696 1197 2 1182 1 1125 NR2P $T=361460 588120 1 0 $X=361460 $Y=582700
X2697 1275 2 1268 1 1141 NR2P $T=373860 699000 1 0 $X=373860 $Y=693580
X2698 1322 2 67 1 1297 NR2P $T=385640 709080 1 180 $X=381920 $Y=708700
X2699 1355 2 1348 1 1362 NR2P $T=391840 598200 0 180 $X=388120 $Y=592780
X2700 1375 2 1367 1 1323 NR2P $T=393080 588120 0 0 $X=393080 $Y=587740
X2701 1391 2 786 1 1241 NR2P $T=402380 658680 0 180 $X=398660 $Y=653260
X2702 1496 2 1477 1 1475 NR2P $T=416020 598200 0 0 $X=416020 $Y=597820
X2703 115 2 114 1 1596 NR2P $T=434000 719160 1 0 $X=434000 $Y=713740
X2704 1646 2 1658 1 1659 NR2P $T=453220 688920 1 180 $X=449500 $Y=688540
X2705 2615 2 2626 1 2634 NR2P $T=685720 598200 1 180 $X=682000 $Y=597820
X2706 2713 2 2628 1 2704 NR2P $T=701840 618360 0 180 $X=698120 $Y=612940
X2707 2782 2 2786 1 2820 NR2P $T=715480 567960 1 180 $X=711760 $Y=567580
X2708 2932 2 2964 1 2965 NR2P $T=734080 628440 1 180 $X=730360 $Y=628060
X2709 2980 2 3018 1 411 NR2P $T=743380 547800 1 0 $X=743380 $Y=542380
X2710 2919 2 3035 1 3150 NR2P $T=761980 658680 0 180 $X=758260 $Y=653260
X2711 3123 2 2965 1 3161 NR2P $T=764460 567960 1 180 $X=760740 $Y=567580
X2712 3105 2 3060 1 3180 NR2P $T=767560 648600 1 180 $X=763840 $Y=648220
X2713 3173 2 3202 1 3215 NR2P $T=770660 688920 1 180 $X=766940 $Y=688540
X2714 3198 2 3233 1 429 NR2P $T=774380 547800 0 180 $X=770660 $Y=542380
X2715 3169 2 3235 1 3270 NR2P $T=778720 598200 1 180 $X=775000 $Y=597820
X2716 430 2 431 1 3278 NR2P $T=781820 547800 0 180 $X=778100 $Y=542380
X2717 3255 2 3286 1 431 NR2P $T=783680 547800 1 180 $X=779960 $Y=547420
X2718 429 2 431 1 435 NR2P $T=781820 547800 1 0 $X=781820 $Y=542380
X2719 3301 2 3254 1 3331 NR2P $T=786780 658680 0 180 $X=783060 $Y=653260
X2720 3228 2 3300 1 3326 NR2P $T=785540 648600 1 0 $X=785540 $Y=643180
X2721 3322 2 3303 1 3334 NR2P $T=789260 668760 0 180 $X=785540 $Y=663340
X2722 3150 2 3301 1 3337 NR2P $T=789880 648600 1 180 $X=786160 $Y=648220
X2723 3336 2 3329 1 3365 NR2P $T=793600 567960 1 180 $X=789880 $Y=567580
X2724 3387 2 3287 1 3404 NR2P $T=799180 588120 0 0 $X=799180 $Y=587740
X2725 3374 2 3393 1 3415 NR2P $T=802900 618360 1 180 $X=799180 $Y=617980
X2726 3314 2 3365 1 3445 NR2P $T=805380 557880 1 180 $X=801660 $Y=557500
X2727 3399 2 3363 1 3447 NR2P $T=807240 588120 0 180 $X=803520 $Y=582700
X2728 3388 2 3214 1 3449 NR2P $T=807240 638520 0 180 $X=803520 $Y=633100
X2729 3447 2 3404 1 3473 NR2P $T=809100 578040 1 180 $X=805380 $Y=577660
X2730 3386 2 3445 1 3439 NR2P $T=806620 557880 0 0 $X=806620 $Y=557500
X2731 3376 2 3417 1 3468 NR2P $T=807860 688920 0 0 $X=807860 $Y=688540
X2732 3415 2 3431 1 3462 NR2P $T=812820 608280 1 180 $X=809100 $Y=607900
X2733 3477 2 3476 1 3466 NR2P $T=811580 709080 1 0 $X=811580 $Y=703660
X2734 3468 2 3485 1 3504 NR2P $T=815920 688920 1 180 $X=812200 $Y=688540
X2735 455 2 453 1 3517 NR2P $T=819640 719160 0 180 $X=815920 $Y=713740
X2736 3510 2 3506 1 3516 NR2P $T=820260 628440 1 0 $X=820260 $Y=623020
X2737 3517 2 3466 1 3505 NR2P $T=820260 699000 0 0 $X=820260 $Y=698620
X2738 3898 2 3945 1 3970 NR2P $T=901480 688920 1 0 $X=901480 $Y=683500
X2739 3969 2 3962 1 3945 NR2P $T=902720 699000 1 0 $X=902720 $Y=693580
X2740 4030 2 4042 1 4023 NR2P $T=916980 688920 1 180 $X=913260 $Y=688540
X2741 4086 2 4106 1 4030 NR2P $T=923800 688920 0 0 $X=923800 $Y=688540
X2742 4201 2 4183 1 4196 NR2P $T=944260 699000 0 0 $X=944260 $Y=698620
X2743 4226 2 602 1 4227 NR2P $T=955420 699000 1 180 $X=951700 $Y=698620
X2744 607 2 604 1 4251 NR2P $T=962240 719160 1 0 $X=962240 $Y=713740
X2745 4329 2 4318 1 4287 NR2P $T=980840 699000 0 0 $X=980840 $Y=698620
X2746 618 2 4318 1 4300 NR2P $T=981460 699000 1 0 $X=981460 $Y=693580
X2747 867 852 1 844 732 842 2 MOAI1 $T=303180 658680 1 180 $X=298840 $Y=658300
X2748 863 851 1 842 850 849 2 MOAI1 $T=304420 638520 1 180 $X=300080 $Y=638140
X2749 851 856 1 842 795 870 2 MOAI1 $T=300700 638520 1 0 $X=300700 $Y=633100
X2750 868 875 1 866 729 864 2 MOAI1 $T=307520 668760 0 180 $X=303180 $Y=663340
X2751 868 871 1 879 817 893 2 MOAI1 $T=303800 648600 1 0 $X=303800 $Y=643180
X2752 872 868 1 883 796 893 2 MOAI1 $T=304420 648600 0 0 $X=304420 $Y=648220
X2753 901 894 1 890 886 882 2 MOAI1 $T=311240 608280 0 180 $X=306900 $Y=602860
X2754 921 867 1 842 888 911 2 MOAI1 $T=315580 658680 1 180 $X=311240 $Y=658300
X2755 868 892 1 937 906 866 2 MOAI1 $T=314960 668760 0 0 $X=314960 $Y=668380
X2756 949 955 1 961 938 968 2 MOAI1 $T=318680 618360 0 0 $X=318680 $Y=617980
X2757 1047 1022 1 1016 823 1012 2 MOAI1 $T=335420 658680 1 180 $X=331080 $Y=658300
X2758 1046 1047 1 1016 791 1066 2 MOAI1 $T=335420 658680 1 0 $X=335420 $Y=653260
X2759 1067 1047 1 1016 998 1086 2 MOAI1 $T=339760 678840 1 0 $X=339760 $Y=673420
X2760 867 1097 1 1106 1111 918 2 MOAI1 $T=345340 618360 1 0 $X=345340 $Y=612940
X2761 1241 1249 1 786 792 1267 2 MOAI1 $T=370140 658680 1 0 $X=370140 $Y=653260
X2762 1185 1301 1 1146 1280 1234 2 MOAI1 $T=381920 638520 0 180 $X=377580 $Y=633100
X2763 1368 1357 1 1363 1347 1342 2 MOAI1 $T=395560 608280 1 180 $X=391220 $Y=607900
X2764 1420 1410 1 1404 1355 1397 2 MOAI1 $T=403000 608280 0 180 $X=398660 $Y=602860
X2765 1433 1428 1 1421 1420 1267 2 MOAI1 $T=407960 648600 1 180 $X=403620 $Y=648220
X2766 1442 1438 1 1430 1418 1427 2 MOAI1 $T=409200 688920 1 180 $X=404860 $Y=688540
X2767 1153 1452 1 1461 1478 1443 2 MOAI1 $T=409200 618360 0 0 $X=409200 $Y=617980
X2768 1241 1538 1 1267 1514 1527 2 MOAI1 $T=429660 648600 1 180 $X=425320 $Y=648220
X2769 107 112 1 113 1557 114 2 MOAI1 $T=429660 719160 1 0 $X=429660 $Y=713740
X2770 125 123 1 121 1598 1335 2 MOAI1 $T=443300 719160 0 180 $X=438960 $Y=713740
X2771 1565 1471 1 1587 1625 1631 2 MOAI1 $T=441440 638520 1 0 $X=441440 $Y=633100
X2772 2644 2657 1 2665 2675 2676 2 MOAI1 $T=687580 578040 1 0 $X=687580 $Y=572620
X2773 2680 2653 1 2735 2751 2743 2 MOAI1 $T=708040 578040 0 180 $X=703700 $Y=572620
X2774 2781 2775 1 2796 2802 2813 2 MOAI1 $T=709900 709080 1 0 $X=709900 $Y=703660
X2775 2658 2772 1 2722 2808 2784 2 MOAI1 $T=717340 618360 1 180 $X=713000 $Y=617980
X2776 2683 2847 1 2815 2814 2829 2 MOAI1 $T=720440 608280 1 180 $X=716100 $Y=607900
X2777 2781 2899 1 2838 2913 2914 2 MOAI1 $T=723540 688920 1 0 $X=723540 $Y=683500
X2778 404 3002 1 405 3001 2996 2 MOAI1 $T=742140 709080 1 180 $X=737800 $Y=708700
X2779 2961 2956 1 3021 3035 2997 2 MOAI1 $T=739040 658680 1 0 $X=739040 $Y=653260
X2780 394 2992 1 3014 3036 3027 2 MOAI1 $T=739040 688920 0 0 $X=739040 $Y=688540
X2781 2959 3006 1 3026 3025 2927 2 MOAI1 $T=740280 598200 1 0 $X=740280 $Y=592780
X2782 407 2979 1 3014 3032 3039 2 MOAI1 $T=740280 709080 1 0 $X=740280 $Y=703660
X2783 407 3043 1 3029 3055 3014 2 MOAI1 $T=744000 688920 0 0 $X=744000 $Y=688540
X2784 2671 3058 1 2678 3034 2984 2 MOAI1 $T=749580 588120 0 180 $X=745240 $Y=582700
X2785 3059 2959 1 2927 3087 3097 2 MOAI1 $T=747100 588120 0 0 $X=747100 $Y=587740
X2786 2910 3042 1 2970 3066 2989 2 MOAI1 $T=752060 618360 0 180 $X=747720 $Y=612940
X2787 3069 2959 1 3083 3092 2927 2 MOAI1 $T=748340 598200 1 0 $X=748340 $Y=592780
X2788 404 3095 1 3014 3088 3081 2 MOAI1 $T=755780 688920 1 180 $X=751440 $Y=688540
X2789 3086 3064 1 3104 3105 3090 2 MOAI1 $T=757640 648600 1 180 $X=753300 $Y=648220
X2790 3130 2918 1 2937 3156 3159 2 MOAI1 $T=758260 618360 0 0 $X=758260 $Y=617980
X2791 2918 3136 1 3127 3147 2937 2 MOAI1 $T=758880 628440 1 0 $X=758880 $Y=623020
X2792 2918 3120 1 3115 3160 2937 2 MOAI1 $T=760120 608280 0 0 $X=760120 $Y=607900
X2793 3108 3139 1 3128 3198 3168 2 MOAI1 $T=763220 547800 0 0 $X=763220 $Y=547420
X2794 3166 3156 1 3178 3203 2943 2 MOAI1 $T=767560 618360 0 0 $X=767560 $Y=617980
X2795 3132 3192 1 3125 3219 3225 2 MOAI1 $T=768800 709080 1 0 $X=768800 $Y=703660
X2796 3238 3132 1 3125 3259 3143 2 MOAI1 $T=775000 719160 1 0 $X=775000 $Y=713740
X2797 3284 3227 1 3288 3430 3296 2 MOAI1 $T=783060 678840 1 0 $X=783060 $Y=673420
X2798 3290 3261 1 3311 3329 3294 2 MOAI1 $T=784300 567960 0 0 $X=784300 $Y=567580
X2799 3369 3243 1 3358 3376 3368 2 MOAI1 $T=799180 699000 0 180 $X=794840 $Y=693580
X2800 536 3871 1 539 542 3921 2 MOAI1 $T=894040 547800 1 0 $X=894040 $Y=542380
X2801 536 3907 1 3928 545 539 2 MOAI1 $T=895900 547800 0 0 $X=895900 $Y=547420
X2802 536 3936 1 3903 3960 3951 2 MOAI1 $T=897760 588120 0 0 $X=897760 $Y=587740
X2803 536 3895 1 3951 552 3955 2 MOAI1 $T=902720 547800 0 0 $X=902720 $Y=547420
X2804 560 4013 1 4038 4045 3951 2 MOAI1 $T=913880 588120 1 0 $X=913880 $Y=582700
X2805 536 4039 1 4053 4058 3951 2 MOAI1 $T=915740 588120 0 0 $X=915740 $Y=587740
X2806 536 4029 1 4060 4063 3951 2 MOAI1 $T=916980 578040 0 0 $X=916980 $Y=577660
X2807 700 1 709 691 2 ND2P $T=265360 658680 1 0 $X=265360 $Y=653260
X2808 708 1 719 715 2 ND2P $T=272180 588120 0 180 $X=268460 $Y=582700
X2809 693 1 714 710 2 ND2P $T=269080 628440 1 0 $X=269080 $Y=623020
X2810 752 1 719 756 2 ND2P $T=279000 578040 0 0 $X=279000 $Y=577660
X2811 784 1 775 779 2 ND2P $T=290160 668760 0 180 $X=286440 $Y=663340
X2812 776 1 719 819 2 ND2P $T=296360 578040 0 0 $X=296360 $Y=577660
X2813 794 1 719 832 2 ND2P $T=297600 588120 1 0 $X=297600 $Y=582700
X2814 846 1 859 847 2 ND2P $T=300700 608280 0 0 $X=300700 $Y=607900
X2815 1107 1 48 46 2 ND2P $T=347200 719160 1 0 $X=347200 $Y=713740
X2816 1122 1 1129 1133 2 ND2P $T=355880 588120 0 0 $X=355880 $Y=587740
X2817 1197 1 1182 1158 2 ND2P $T=364560 588120 1 180 $X=360840 $Y=587740
X2818 1225 1 1199 1144 2 ND2P $T=367660 699000 0 0 $X=367660 $Y=698620
X2819 1275 1 1268 1181 2 ND2P $T=378200 699000 1 0 $X=378200 $Y=693580
X2820 1324 1 1323 1302 2 ND2P $T=386260 578040 1 180 $X=382540 $Y=577660
X2821 1441 1 1426 1379 2 ND2P $T=407340 678840 0 0 $X=407340 $Y=678460
X2822 1544 1 1581 1543 2 ND2P $T=434620 598200 0 0 $X=434620 $Y=597820
X2823 1562 1 1585 1487 2 ND2P $T=435240 678840 0 0 $X=435240 $Y=678460
X2824 1632 1 1636 1602 2 ND2P $T=445780 678840 1 0 $X=445780 $Y=673420
X2825 2648 1 2638 2654 2 ND2P $T=688200 608280 1 0 $X=688200 $Y=602860
X2826 378 1 375 2817 2 ND2P $T=714860 547800 0 180 $X=711140 $Y=542380
X2827 2881 1 2862 2871 2 ND2P $T=723540 598200 0 0 $X=723540 $Y=597820
X2828 3283 1 3280 3314 2 ND2P $T=790500 557880 1 180 $X=786780 $Y=557500
X2829 3321 1 3331 3309 2 ND2P $T=787400 658680 0 0 $X=787400 $Y=658300
X2830 3337 1 3321 3348 2 ND2P $T=795460 648600 1 180 $X=791740 $Y=648220
X2831 3327 1 3236 3345 2 ND2P $T=795460 668760 1 180 $X=791740 $Y=668380
X2832 3383 1 3295 3412 2 ND2P $T=798560 618360 1 0 $X=798560 $Y=612940
X2833 3399 1 3363 3402 2 ND2P $T=803520 588120 0 180 $X=799800 $Y=582700
X2834 451 1 449 3477 2 ND2P $T=809100 719160 0 180 $X=805380 $Y=713740
X2835 3443 1 3461 3446 2 ND2P $T=807240 598200 0 0 $X=807240 $Y=597820
X2836 455 1 453 3464 2 ND2P $T=815300 719160 0 180 $X=811580 $Y=713740
X2837 3462 1 3461 3491 2 ND2P $T=816540 598200 0 0 $X=816540 $Y=597820
X2838 3530 1 3461 3535 2 ND2P $T=821500 608280 1 0 $X=821500 $Y=602860
X2839 514 1 515 3742 2 ND2P $T=871720 719160 1 0 $X=871720 $Y=713740
X2840 4023 1 3983 4102 2 ND2P $T=918220 688920 1 0 $X=918220 $Y=683500
X2841 4287 1 4264 4308 2 ND2P $T=974640 699000 0 180 $X=970920 $Y=693580
X2842 791 778 796 1 2 741 MAO222 $T=292640 648600 0 180 $X=287680 $Y=643180
X2843 751 746 733 1 2 762 MAO222 $T=293260 618360 1 180 $X=288300 $Y=617980
X2844 888 877 907 1 2 763 MAO222 $T=309380 678840 1 180 $X=304420 $Y=678460
X2845 906 904 896 1 2 814 MAO222 $T=308760 678840 1 0 $X=308760 $Y=673420
X2846 1163 1169 1190 1 2 1108 MAO222 $T=362080 598200 1 180 $X=357120 $Y=597820
X2847 1253 1261 1235 1 2 1251 MAO222 $T=375720 598200 1 180 $X=370760 $Y=597820
X2848 1372 1384 1398 1 2 1368 MAO222 $T=399280 638520 0 180 $X=394320 $Y=633100
X2849 100 1503 1469 1 2 1442 MAO222 $T=417260 699000 1 0 $X=417260 $Y=693580
X2850 117 1583 1557 1 2 1589 MAO222 $T=435240 688920 0 0 $X=435240 $Y=688540
X2851 126 1617 1596 1 2 1626 MAO222 $T=442060 709080 1 0 $X=442060 $Y=703660
X2852 2814 2810 2790 1 2 2860 MAO222 $T=716100 557880 0 0 $X=716100 $Y=557500
X2853 2857 2849 2720 1 2 2890 MAO222 $T=719820 588120 0 0 $X=719820 $Y=587740
X2854 2966 2981 2934 1 2 3037 MAO222 $T=739660 557880 0 0 $X=739660 $Y=557500
X2855 3047 412 2973 1 2 3064 MAO222 $T=743380 678840 1 0 $X=743380 $Y=673420
X2856 3034 3077 2978 1 2 3108 MAO222 $T=750820 567960 1 0 $X=750820 $Y=562540
X2857 3036 3153 3122 1 2 3187 MAO222 $T=762600 668760 0 0 $X=762600 $Y=668380
X2858 3148 3054 3025 1 2 3184 MAO222 $T=763220 557880 0 0 $X=763220 $Y=557500
X2859 3161 3154 3052 1 2 3207 MAO222 $T=765700 567960 0 0 $X=765700 $Y=567580
X2860 3138 3209 3055 1 2 3232 MAO222 $T=769420 678840 1 0 $X=769420 $Y=673420
X2861 3184 3211 3176 1 2 3255 MAO222 $T=772520 557880 1 0 $X=772520 $Y=552460
X2862 3032 3272 3258 1 2 3292 MAO222 $T=778720 709080 1 0 $X=778720 $Y=703660
X2863 3245 3269 3092 1 2 3312 MAO222 $T=779340 588120 1 0 $X=779340 $Y=582700
X2864 433 436 434 1 2 3310 MAO222 $T=781820 719160 1 0 $X=781820 $Y=713740
X2865 3253 3165 3256 1 2 3327 MAO222 $T=784300 678840 0 0 $X=784300 $Y=678460
X2866 3160 3299 3212 1 2 3347 MAO222 $T=785540 608280 0 0 $X=785540 $Y=607900
X2867 529 525 530 1 2 3844 MAO222 $T=890940 719160 0 180 $X=885980 $Y=713740
X2868 582 4143 578 1 2 4173 MAO222 $T=933720 709080 0 0 $X=933720 $Y=708700
X2869 4198 4319 4336 1 2 625 MAO222 $T=986420 598200 1 0 $X=986420 $Y=592780
X2870 709 687 2 689 723 1 678 FA1 $T=272800 658680 1 180 $X=257300 $Y=658300
X2871 723 729 2 732 759 1 697 FA1 $T=283960 668760 0 180 $X=268460 $Y=663340
X2872 775 763 2 765 802 1 700 FA1 $T=294500 678840 1 180 $X=279000 $Y=678460
X2873 695 786 2 799 850 1 702 FA1 $T=279620 638520 0 0 $X=279620 $Y=638140
X2874 733 895 2 897 848 1 787 FA1 $T=298840 618360 0 0 $X=298840 $Y=617980
X2875 747 799 2 874 878 1 848 FA1 $T=315580 628440 1 180 $X=300080 $Y=628060
X2876 751 919 2 929 936 1 894 FA1 $T=303800 628440 1 0 $X=303800 $Y=623020
X2877 901 1010 2 1045 1019 1 1069 FA1 $T=324880 618360 0 0 $X=324880 $Y=617980
X2878 899 1036 2 1064 1069 1 1072 FA1 $T=329220 618360 1 0 $X=329220 $Y=612940
X2879 1036 1090 2 1077 1054 1 1089 FA1 $T=334800 628440 1 0 $X=334800 $Y=623020
X2880 1129 1108 2 1102 1115 1 1033 FA1 $T=358360 598200 0 180 $X=342860 $Y=592780
X2881 1182 1203 2 1205 1251 1 1122 FA1 $T=375100 598200 0 180 $X=359600 $Y=592780
X2882 1268 1288 2 65 1331 1 1199 FA1 $T=388120 699000 1 180 $X=372620 $Y=698620
X2883 1534 1492 2 1478 1519 1 1466 FA1 $T=427800 608280 1 180 $X=412300 $Y=607900
X2884 1548 1514 2 1506 1518 1 1493 FA1 $T=432760 618360 1 180 $X=417260 $Y=617980
X2885 2723 2708 2 2721 2763 1 2692 FA1 $T=710520 678840 1 180 $X=695020 $Y=678460
X2886 2788 2723 2 2725 2769 1 2693 FA1 $T=711140 668760 0 180 $X=695640 $Y=663340
X2887 2956 388 2 384 2836 1 2823 FA1 $T=730360 668760 1 180 $X=714860 $Y=668380
X2888 2985 2897 2 2891 2873 1 2835 FA1 $T=735320 648600 1 180 $X=719820 $Y=648220
X2889 3013 2938 2 2806 2923 1 2873 FA1 $T=740900 648600 0 180 $X=725400 $Y=643180
X2890 2971 2954 2 2878 2993 1 3075 FA1 $T=734700 608280 0 0 $X=734700 $Y=607900
X2891 3086 3022 2 3000 2990 1 2988 FA1 $T=752060 668760 0 180 $X=736560 $Y=663340
X2892 3091 2707 2 2785 3030 1 3201 FA1 $T=753300 638520 0 0 $X=753300 $Y=638140
X2893 3303 3187 2 3065 3140 1 3155 FA1 $T=778100 668760 0 180 $X=762600 $Y=663340
X2894 3163 3213 2 3066 3075 1 3281 FA1 $T=764460 618360 1 0 $X=764460 $Y=612940
X2895 3196 3244 2 3087 3146 1 3290 FA1 $T=769420 578040 1 0 $X=769420 $Y=572620
X2896 3214 3013 2 3201 3208 1 3333 FA1 $T=771280 638520 0 0 $X=771280 $Y=638140
X2897 3236 3232 2 3131 3218 1 3322 FA1 $T=774380 668760 0 0 $X=774380 $Y=668380
X2898 3287 3347 2 3276 3163 1 3383 FA1 $T=782440 618360 1 0 $X=782440 $Y=612940
X2899 3295 3340 2 3203 3281 1 3393 FA1 $T=783680 618360 0 0 $X=783680 $Y=617980
X2900 3529 3569 2 474 2323 1 3619 FA1 $T=822740 588120 1 0 $X=822740 $Y=582700
X2901 3539 3581 2 472 2278 1 3583 FA1 $T=824600 598200 1 0 $X=824600 $Y=592780
X2902 3552 3575 2 3521 2254 1 3636 FA1 $T=828940 598200 0 0 $X=828940 $Y=597820
X2903 3565 3620 2 483 2307 1 485 FA1 $T=832040 567960 1 0 $X=832040 $Y=562540
X2904 3962 567 2 568 556 1 4043 FA1 $T=907680 709080 0 0 $X=907680 $Y=708700
X2905 4154 4173 2 591 4186 1 4201 FA1 $T=934340 709080 1 0 $X=934340 $Y=703660
X2906 4183 598 2 4217 592 1 4226 FA1 $T=941780 709080 0 0 $X=941780 $Y=708700
X2907 684 704 2 1 717 OR2 $T=267220 608280 1 0 $X=267220 $Y=602860
X2908 795 817 2 1 797 OR2 $T=296360 628440 1 180 $X=293880 $Y=628060
X2909 972 958 2 1 820 OR2 $T=321780 678840 1 180 $X=319300 $Y=678460
X2910 1040 1038 2 1 43 OR2 $T=344100 547800 0 0 $X=344100 $Y=547420
X2911 1136 1150 2 1 961 OR2 $T=354640 628440 1 0 $X=354640 $Y=623020
X2912 1334 1340 2 1 1317 OR2 $T=388740 688920 1 180 $X=386260 $Y=688540
X2913 75 70 2 1 1385 OR2 $T=393700 719160 1 0 $X=393700 $Y=713740
X2914 1460 1466 2 1 1508 OR2 $T=420360 598200 0 0 $X=420360 $Y=597820
X2915 1534 1493 2 1 1521 OR2 $T=426560 608280 0 180 $X=424080 $Y=602860
X2916 1550 1561 2 1 1574 OR2 $T=432760 618360 0 0 $X=432760 $Y=617980
X2917 1547 1589 2 1 1599 OR2 $T=438340 688920 1 0 $X=438340 $Y=683500
X2918 1601 1605 2 1 1642 OR2 $T=446400 638520 1 0 $X=446400 $Y=633100
X2919 1678 1664 2 1 1675 OR2 $T=456320 709080 1 0 $X=456320 $Y=703660
X2920 1744 1727 2 1 1769 OR2 $T=469960 608280 0 0 $X=469960 $Y=607900
X2921 2691 2686 2 1 362 OR2 $T=696260 547800 1 180 $X=693780 $Y=547420
X2922 2700 2711 2 1 2655 OR2 $T=700600 567960 0 180 $X=698120 $Y=562540
X2923 2706 2717 2 1 2746 OR2 $T=701840 557880 1 0 $X=701840 $Y=552460
X2924 2751 2747 2 1 2742 OR2 $T=706180 567960 0 180 $X=703700 $Y=562540
X2925 2699 2803 2 1 2827 OR2 $T=712380 588120 1 0 $X=712380 $Y=582700
X2926 2818 2768 2 1 383 OR2 $T=715480 547800 0 0 $X=715480 $Y=547420
X2927 2866 2739 2 1 2881 OR2 $T=721060 598200 0 0 $X=721060 $Y=597820
X2928 2735 2825 2 1 2901 OR2 $T=727260 588120 1 180 $X=724780 $Y=587740
X2929 3207 3239 2 1 3248 OR2 $T=774380 567960 0 0 $X=774380 $Y=567580
X2930 3150 3158 2 1 3254 OR2 $T=774380 658680 1 0 $X=774380 $Y=653260
X2931 3228 3150 2 1 3343 OR2 $T=789880 648600 1 0 $X=789880 $Y=643180
X2932 3292 3242 2 1 3378 OR2 $T=794220 688920 0 0 $X=794220 $Y=688540
X2933 3447 3439 2 1 3423 OR2 $T=806620 567960 1 180 $X=804140 $Y=567580
X2934 3442 3444 2 1 3482 OR2 $T=808480 678840 0 0 $X=808480 $Y=678460
X2935 3445 3386 2 1 3500 OR2 $T=812200 557880 0 0 $X=812200 $Y=557500
X2936 3451 3508 2 1 3515 OR2 $T=817160 668760 0 0 $X=817160 $Y=668380
X2937 3487 3449 2 1 3522 OR2 $T=818400 618360 1 0 $X=818400 $Y=612940
X2938 3555 3546 2 1 3545 OR2 $T=829560 618360 0 180 $X=827080 $Y=612940
X2939 3648 3658 2 1 3680 OR2 $T=848780 618360 1 0 $X=848780 $Y=612940
X2940 522 3788 2 1 3771 OR2 $T=877300 709080 1 180 $X=874820 $Y=708700
X2941 3840 3844 2 1 3785 OR2 $T=884120 699000 0 0 $X=884120 $Y=698620
X2942 3855 3753 2 1 3896 OR2 $T=890320 588120 0 0 $X=890320 $Y=587740
X2943 3979 3831 2 1 3991 OR2 $T=906440 598200 0 0 $X=906440 $Y=597820
X2944 4025 3992 2 1 4003 OR2 $T=913260 557880 1 180 $X=910780 $Y=557500
X2945 4057 4036 2 1 4019 OR2 $T=916980 648600 1 180 $X=914500 $Y=648220
X2946 4218 4227 2 1 4241 OR2 $T=954180 678840 0 0 $X=954180 $Y=678460
X2947 860 811 2 873 1 910 AOI12HS $T=307520 588120 0 0 $X=307520 $Y=587740
X2948 18 21 2 898 1 933 AOI12HS $T=316820 547800 0 180 $X=312480 $Y=542380
X2949 43 32 2 1063 1 1081 AOI12HS $T=344720 547800 0 180 $X=340380 $Y=542380
X2950 1035 959 2 922 1 1075 AOI12HS $T=344100 578040 0 0 $X=344100 $Y=577660
X2951 1099 1062 2 1060 1 1130 AOI12HS $T=347200 699000 1 0 $X=347200 $Y=693580
X2952 1135 1145 2 1151 1 28 AOI12HS $T=352780 557880 1 0 $X=352780 $Y=552460
X2953 1135 1145 2 1151 1 952 AOI12HS $T=354020 547800 0 0 $X=354020 $Y=547420
X2954 1156 1152 2 1120 1 1142 AOI12HS $T=358360 567960 0 180 $X=354020 $Y=562540
X2955 1166 1035 2 1184 1 1159 AOI12HS $T=358980 578040 0 0 $X=358980 $Y=577660
X2956 1215 1153 2 1188 1 1176 AOI12HS $T=367040 618360 0 180 $X=362700 $Y=612940
X2957 1212 1229 2 1178 1 1237 AOI12HS $T=370760 567960 1 180 $X=366420 $Y=567580
X2958 1226 1229 2 1245 1 1232 AOI12HS $T=367660 557880 0 0 $X=367660 $Y=557500
X2959 1172 1229 2 1156 1 1254 AOI12HS $T=372000 567960 0 180 $X=367660 $Y=562540
X2960 1260 1099 2 1242 1 1214 AOI12HS $T=373240 688920 1 180 $X=368900 $Y=688540
X2961 62 1250 2 59 1 1167 AOI12HS $T=375720 547800 0 180 $X=371380 $Y=542380
X2962 1339 1353 2 976 1 1274 AOI12HS $T=389360 618360 1 180 $X=385020 $Y=617980
X2963 1361 1354 2 1323 1 1373 AOI12HS $T=398040 578040 1 180 $X=393700 $Y=577660
X2964 1487 1467 2 1441 1 1437 AOI12HS $T=417260 678840 0 180 $X=412920 $Y=673420
X2965 1600 1610 2 1620 1 1604 AOI12HS $T=440200 618360 1 0 $X=440200 $Y=612940
X2966 1690 1675 2 1670 1 1653 AOI12HS $T=458180 699000 1 180 $X=453840 $Y=698620
X2967 1738 1730 2 1709 1 1737 AOI12HS $T=471200 547800 1 180 $X=466860 $Y=547420
X2968 1767 1769 2 1782 1 1786 AOI12HS $T=473060 608280 0 0 $X=473060 $Y=607900
X2969 1772 1783 2 1738 1 1792 AOI12HS $T=474300 557880 1 0 $X=474300 $Y=552460
X2970 1795 1783 2 1753 1 1762 AOI12HS $T=479260 557880 1 180 $X=474920 $Y=557500
X2971 1774 1785 2 1768 1 1746 AOI12HS $T=475540 578040 0 0 $X=475540 $Y=577660
X2972 1799 1783 2 1829 1 1841 AOI12HS $T=481120 578040 1 0 $X=481120 $Y=572620
X2973 2662 2704 2 2663 1 2696 AOI12HS $T=700600 608280 1 180 $X=696260 $Y=607900
X2974 2930 394 2 2948 1 2753 AOI12HS $T=728500 688920 1 0 $X=728500 $Y=683500
X2975 3381 3385 2 3398 1 3357 AOI12HS $T=796700 557880 1 0 $X=796700 $Y=552460
X2976 3486 3385 2 3500 1 3467 AOI12HS $T=812820 567960 1 0 $X=812820 $Y=562540
X2977 3490 3420 2 3487 1 3511 AOI12HS $T=814060 618360 1 0 $X=814060 $Y=612940
X2978 3551 3544 2 3537 1 3554 AOI12HS $T=828940 709080 0 180 $X=824600 $Y=703660
X2979 3505 3544 2 3499 1 3550 AOI12HS $T=827700 699000 1 0 $X=827700 $Y=693580
X2980 3593 3591 2 3576 1 3585 AOI12HS $T=837620 688920 0 180 $X=833280 $Y=683500
X2981 3598 3545 2 3587 1 3612 AOI12HS $T=840100 618360 0 180 $X=835760 $Y=612940
X2982 3622 3591 2 3605 1 3613 AOI12HS $T=842580 678840 1 180 $X=838240 $Y=678460
X2983 3605 3617 2 3629 1 3639 AOI12HS $T=840100 699000 1 0 $X=840100 $Y=693580
X2984 3645 3660 2 3670 1 3678 AOI12HS $T=846920 557880 1 0 $X=846920 $Y=552460
X2985 3654 3591 2 3642 1 3676 AOI12HS $T=846920 678840 0 0 $X=846920 $Y=678460
X2986 3665 3685 2 3677 1 3688 AOI12HS $T=855600 578040 0 180 $X=851260 $Y=572620
X2987 3771 3742 2 3749 1 3752 AOI12HS $T=872960 699000 1 180 $X=868620 $Y=698620
X2988 3768 3769 2 3750 1 3756 AOI12HS $T=874200 557880 0 180 $X=869860 $Y=552460
X2989 3776 518 2 3768 1 3803 AOI12HS $T=874200 547800 0 0 $X=874200 $Y=547420
X2990 3781 3773 2 3797 1 3789 AOI12HS $T=874820 648600 0 0 $X=874820 $Y=648220
X2991 3795 518 2 3813 1 3825 AOI12HS $T=877300 557880 1 0 $X=877300 $Y=552460
X2992 3773 3811 2 3818 1 3809 AOI12HS $T=879160 648600 0 0 $X=879160 $Y=648220
X2993 3837 3852 2 3858 1 3847 AOI12HS $T=884740 638520 0 0 $X=884740 $Y=638140
X2994 3849 3663 2 3861 1 3864 AOI12HS $T=885360 648600 1 0 $X=885360 $Y=643180
X2995 3881 3862 2 3857 1 3866 AOI12HS $T=890320 688920 1 180 $X=885980 $Y=688540
X2996 3867 3846 2 3868 1 3908 AOI12HS $T=894660 578040 1 180 $X=890320 $Y=577660
X2997 3885 3852 2 3909 1 3914 AOI12HS $T=893420 648600 1 0 $X=893420 $Y=643180
X2998 3909 3932 2 3941 1 3880 AOI12HS $T=897140 648600 0 0 $X=897140 $Y=648220
X2999 3922 3867 2 3946 1 3938 AOI12HS $T=897760 578040 0 0 $X=897760 $Y=577660
X3000 3891 3852 2 3947 1 3913 AOI12HS $T=897760 638520 1 0 $X=897760 $Y=633100
X3001 3950 3917 2 3973 1 3978 AOI12HS $T=902720 588120 1 0 $X=902720 $Y=582700
X3002 3896 3917 2 3974 1 3995 AOI12HS $T=903960 598200 1 0 $X=903960 $Y=592780
X3003 3862 3970 2 3983 1 3954 AOI12HS $T=903960 678840 0 0 $X=903960 $Y=678460
X3004 3971 3917 2 3990 1 4004 AOI12HS $T=905200 578040 0 0 $X=905200 $Y=577660
X3005 3974 3991 2 4005 1 3981 AOI12HS $T=907060 588120 0 0 $X=907060 $Y=587740
X3006 3998 4003 2 4012 1 3989 AOI12HS $T=908920 567960 1 0 $X=908920 $Y=562540
X3007 4019 4018 2 4055 1 4032 AOI12HS $T=915120 638520 0 0 $X=915120 $Y=638140
X3008 4040 547 2 4059 1 569 AOI12HS $T=916360 547800 1 0 $X=916360 $Y=542380
X3009 4097 4103 2 4114 1 4123 AOI12HS $T=923800 578040 0 0 $X=923800 $Y=577660
X3010 4119 4113 2 4138 1 4088 AOI12HS $T=927520 557880 0 0 $X=927520 $Y=557500
X3011 4136 4103 2 4111 1 4148 AOI12HS $T=935580 567960 1 180 $X=931240 $Y=567580
X3012 4105 4103 2 4119 1 4139 AOI12HS $T=937440 578040 0 180 $X=933100 $Y=572620
X3013 4150 4124 2 4160 1 4149 AOI12HS $T=933100 628440 0 0 $X=933100 $Y=628060
X3014 4124 4159 2 4161 1 4095 AOI12HS $T=933100 638520 0 0 $X=933100 $Y=638140
X3015 4180 4162 2 4193 1 4192 AOI12HS $T=941160 688920 0 0 $X=941160 $Y=688540
X3016 4200 4129 2 4210 1 4209 AOI12HS $T=945500 678840 0 0 $X=945500 $Y=678460
X3017 4249 4129 2 4264 1 4258 AOI12HS $T=959760 688920 1 0 $X=959760 $Y=683500
X3018 695 697 706 2 1 XOR2HS $T=263500 648600 0 0 $X=263500 $Y=648220
X3019 726 730 740 2 1 XOR2HS $T=272800 578040 1 0 $X=272800 $Y=572620
X3020 791 796 773 2 1 XOR2HS $T=293260 658680 0 180 $X=287680 $Y=653260
X3021 810 814 829 2 1 XOR2HS $T=293260 688920 0 0 $X=293260 $Y=688540
X3022 828 837 845 2 1 XOR2HS $T=296360 678840 1 0 $X=296360 $Y=673420
X3023 838 910 924 2 1 XOR2HS $T=312480 588120 0 0 $X=312480 $Y=587740
X3024 939 932 856 2 1 XOR2HS $T=318680 648600 0 180 $X=313100 $Y=643180
X3025 939 963 876 2 1 XOR2HS $T=323020 668760 0 180 $X=317440 $Y=663340
X3026 939 974 934 2 1 XOR2HS $T=324880 648600 0 180 $X=319300 $Y=643180
X3027 939 977 852 2 1 XOR2HS $T=325500 658680 1 180 $X=319920 $Y=658300
X3028 955 949 981 2 1 XOR2HS $T=322400 628440 1 0 $X=322400 $Y=623020
X3029 871 977 892 2 1 XOR2HS $T=327980 668760 1 180 $X=322400 $Y=668380
X3030 983 989 891 2 1 XOR2HS $T=329220 638520 0 180 $X=323640 $Y=633100
X3031 1017 1061 927 2 1 XOR2HS $T=341000 628440 1 180 $X=335420 $Y=628060
X3032 1053 1075 1056 2 1 XOR2HS $T=344100 578040 1 180 $X=338520 $Y=577660
X3033 1049 1055 1000 2 1 XOR2HS $T=344100 668760 1 180 $X=338520 $Y=668380
X3034 1092 1001 1058 2 1 XOR2HS $T=345960 668760 0 180 $X=340380 $Y=663340
X3035 983 1109 946 2 1 XOR2HS $T=349680 628440 1 180 $X=344100 $Y=628060
X3036 1023 952 1127 2 1 XOR2HS $T=347820 547800 0 0 $X=347820 $Y=547420
X3037 1118 1130 1140 2 1 XOR2HS $T=350300 688920 0 0 $X=350300 $Y=688540
X3038 1092 1109 1067 2 1 XOR2HS $T=357740 678840 0 180 $X=352160 $Y=673420
X3039 1018 50 1160 2 1 XOR2HS $T=363320 658680 0 180 $X=357740 $Y=653260
X3040 1209 914 1187 2 1 XOR2HS $T=366420 678840 1 180 $X=360840 $Y=678460
X3041 1176 1190 1206 2 1 XOR2HS $T=361460 608280 1 0 $X=361460 $Y=602860
X3042 1209 977 1191 2 1 XOR2HS $T=367040 668760 0 180 $X=361460 $Y=663340
X3043 983 1131 1215 2 1 XOR2HS $T=362700 628440 1 0 $X=362700 $Y=623020
X3044 1209 974 1249 2 1 XOR2HS $T=367040 658680 0 0 $X=367040 $Y=658300
X3045 1209 989 1244 2 1 XOR2HS $T=367040 668760 1 0 $X=367040 $Y=663340
X3046 1209 932 1216 2 1 XOR2HS $T=367040 678840 0 0 $X=367040 $Y=678460
X3047 1236 1223 1257 2 1 XOR2HS $T=368900 628440 1 0 $X=368900 $Y=623020
X3048 1147 1189 1264 2 1 XOR2HS $T=370760 638520 0 0 $X=370760 $Y=638140
X3049 1209 963 1183 2 1 XOR2HS $T=378820 668760 0 180 $X=373240 $Y=663340
X3050 1253 1293 1290 2 1 XOR2HS $T=377580 598200 1 0 $X=377580 $Y=592780
X3051 1235 1261 1293 2 1 XOR2HS $T=377580 598200 0 0 $X=377580 $Y=597820
X3052 1306 1001 1269 2 1 XOR2HS $T=388740 668760 0 180 $X=383160 $Y=663340
X3053 1280 1314 1342 2 1 XOR2HS $T=384400 608280 0 0 $X=384400 $Y=607900
X3054 1321 1332 1357 2 1 XOR2HS $T=386880 638520 1 0 $X=386880 $Y=633100
X3055 1306 50 1337 2 1 XOR2HS $T=393700 658680 1 180 $X=388120 $Y=658300
X3056 1357 1368 1356 2 1 XOR2HS $T=394940 608280 0 180 $X=389360 $Y=602860
X3057 1349 1373 1346 2 1 XOR2HS $T=396180 578040 0 180 $X=390600 $Y=572620
X3058 1313 1017 1202 2 1 XOR2HS $T=396800 628440 1 180 $X=391220 $Y=628060
X3059 1341 71 1380 2 1 XOR2HS $T=391840 709080 1 0 $X=391840 $Y=703660
X3060 1306 1109 1369 2 1 XOR2HS $T=393700 658680 0 0 $X=393700 $Y=658300
X3061 1361 1388 1413 2 1 XOR2HS $T=398040 578040 0 0 $X=398040 $Y=577660
X3062 1384 1423 1404 2 1 XOR2HS $T=405480 628440 1 180 $X=399900 $Y=628060
X3063 1410 1420 1440 2 1 XOR2HS $T=404240 608280 0 0 $X=404240 $Y=607900
X3064 1429 1437 1449 2 1 XOR2HS $T=405480 678840 1 0 $X=405480 $Y=673420
X3065 1408 1315 1452 2 1 XOR2HS $T=406100 628440 1 0 $X=406100 $Y=623020
X3066 1223 1344 1474 2 1 XOR2HS $T=410440 638520 1 0 $X=410440 $Y=633100
X3067 1306 1155 1428 2 1 XOR2HS $T=411060 658680 1 0 $X=411060 $Y=653260
X3068 1465 1476 1486 2 1 XOR2HS $T=412920 688920 1 0 $X=412920 $Y=683500
X3069 1131 1453 1504 2 1 XOR2HS $T=416640 658680 1 0 $X=416640 $Y=653260
X3070 1453 1472 1513 2 1 XOR2HS $T=418500 648600 1 0 $X=418500 $Y=643180
X3071 1503 1507 1532 2 1 XOR2HS $T=422840 699000 0 0 $X=422840 $Y=698620
X3072 1487 1522 1546 2 1 XOR2HS $T=425940 678840 1 0 $X=425940 $Y=673420
X3073 105 1516 1567 2 1 XOR2HS $T=429660 699000 1 0 $X=429660 $Y=693580
X3074 1566 1223 1538 2 1 XOR2HS $T=436480 638520 1 180 $X=430900 $Y=638140
X3075 1583 117 1607 2 1 XOR2HS $T=437100 699000 1 0 $X=437100 $Y=693580
X3076 1566 1339 1565 2 1 XOR2HS $T=438340 628440 0 0 $X=438340 $Y=628060
X3077 1581 1569 1619 2 1 XOR2HS $T=440200 598200 0 0 $X=440200 $Y=597820
X3078 1617 1596 1630 2 1 XOR2HS $T=441440 699000 0 0 $X=441440 $Y=698620
X3079 1604 1612 1633 2 1 XOR2HS $T=442680 608280 1 0 $X=442680 $Y=602860
X3080 126 1630 1649 2 1 XOR2HS $T=447020 699000 0 0 $X=447020 $Y=698620
X3081 1636 1629 1663 2 1 XOR2HS $T=450120 678840 1 0 $X=450120 $Y=673420
X3082 1642 1657 1654 2 1 XOR2HS $T=450740 628440 1 0 $X=450740 $Y=623020
X3083 1566 1189 1608 2 1 XOR2HS $T=458800 638520 1 180 $X=453220 $Y=638140
X3084 1653 1683 1682 2 1 XOR2HS $T=456940 688920 1 0 $X=456940 $Y=683500
X3085 141 1721 1726 2 1 XOR2HS $T=464380 709080 1 0 $X=464380 $Y=703660
X3086 1711 1762 1771 2 1 XOR2HS $T=471200 547800 0 0 $X=471200 $Y=547420
X3087 1786 1796 1807 2 1 XOR2HS $T=477400 598200 0 0 $X=477400 $Y=597820
X3088 1798 1792 1818 2 1 XOR2HS $T=478640 557880 1 0 $X=478640 $Y=552460
X3089 1820 1784 1849 2 1 XOR2HS $T=482980 598200 1 0 $X=482980 $Y=592780
X3090 1763 1841 1857 2 1 XOR2HS $T=486080 578040 1 0 $X=486080 $Y=572620
X3091 2615 2626 2622 2 1 XOR2HS $T=683860 598200 0 180 $X=678280 $Y=592780
X3092 2655 2650 356 2 1 XOR2HS $T=689440 567960 0 180 $X=683860 $Y=562540
X3093 2626 2642 2653 2 1 XOR2HS $T=684480 588120 1 0 $X=684480 $Y=582700
X3094 2662 2637 2644 2 1 XOR2HS $T=690680 578040 1 180 $X=685100 $Y=577660
X3095 2639 2628 2658 2 1 XOR2HS $T=685100 618360 0 0 $X=685100 $Y=617980
X3096 2628 2642 2677 2 1 XOR2HS $T=688820 618360 1 0 $X=688820 $Y=612940
X3097 2673 2642 2684 2 1 XOR2HS $T=691300 598200 1 0 $X=691300 $Y=592780
X3098 2637 2727 2698 2 1 XOR2HS $T=703080 578040 1 180 $X=697500 $Y=577660
X3099 2664 2732 364 2 1 XOR2HS $T=704320 547800 0 180 $X=698740 $Y=542380
X3100 2663 2662 2712 2 1 XOR2HS $T=699980 588120 0 0 $X=699980 $Y=587740
X3101 2726 2693 2750 2 1 XOR2HS $T=701220 658680 0 0 $X=701220 $Y=658300
X3102 2727 2673 2761 2 1 XOR2HS $T=703700 598200 1 0 $X=703700 $Y=592780
X3103 2733 370 2770 2 1 XOR2HS $T=704320 699000 0 0 $X=704320 $Y=698620
X3104 2744 2754 2771 2 1 XOR2HS $T=704940 557880 1 0 $X=704940 $Y=552460
X3105 2727 2631 2772 2 1 XOR2HS $T=704940 628440 1 0 $X=704940 $Y=623020
X3106 2651 2727 2774 2 1 XOR2HS $T=705560 598200 0 0 $X=705560 $Y=597820
X3107 2765 2651 2794 2 1 XOR2HS $T=708660 608280 1 0 $X=708660 $Y=602860
X3108 2637 2719 2787 2 1 XOR2HS $T=710520 578040 0 0 $X=710520 $Y=577660
X3109 2645 2663 2803 2 1 XOR2HS $T=711760 598200 1 0 $X=711760 $Y=592780
X3110 2820 2834 2854 2 1 XOR2HS $T=715480 567960 1 0 $X=715480 $Y=562540
X3111 2819 2835 2856 2 1 XOR2HS $T=715480 658680 1 0 $X=715480 $Y=653260
X3112 2861 2855 2834 2 1 XOR2HS $T=721680 567960 1 180 $X=716100 $Y=567580
X3113 366 374 387 2 1 XOR2HS $T=716100 719160 1 0 $X=716100 $Y=713740
X3114 2871 2865 2846 2 1 XOR2HS $T=722920 557880 0 180 $X=717340 $Y=552460
X3115 2837 2645 2870 2 1 XOR2HS $T=717960 608280 1 0 $X=717960 $Y=602860
X3116 2846 2854 2876 2 1 XOR2HS $T=719200 547800 0 0 $X=719200 $Y=547420
X3117 2718 2630 2886 2 1 XOR2HS $T=720440 608280 0 0 $X=720440 $Y=607900
X3118 2830 391 2858 2 1 XOR2HS $T=727260 699000 1 180 $X=721680 $Y=698620
X3119 2906 2792 2922 2 1 XOR2HS $T=732220 578040 1 180 $X=726640 $Y=577660
X3120 2830 400 2899 2 1 XOR2HS $T=732840 699000 1 180 $X=727260 $Y=698620
X3121 2900 373 2930 2 1 XOR2HS $T=733460 688920 1 180 $X=727880 $Y=688540
X3122 371 2921 401 2 1 XOR2HS $T=727880 709080 0 0 $X=727880 $Y=708700
X3123 2943 2630 2962 2 1 XOR2HS $T=730980 608280 1 0 $X=730980 $Y=602860
X3124 2900 370 2979 2 1 XOR2HS $T=732220 709080 1 0 $X=732220 $Y=703660
X3125 2951 2939 2944 2 1 XOR2HS $T=733460 658680 0 0 $X=733460 $Y=658300
X3126 2900 376 2968 2 1 XOR2HS $T=733460 688920 1 0 $X=733460 $Y=683500
X3127 2900 389 2991 2 1 XOR2HS $T=733460 688920 0 0 $X=733460 $Y=688540
X3128 2900 400 2992 2 1 XOR2HS $T=733460 699000 0 0 $X=733460 $Y=698620
X3129 2906 2715 2974 2 1 XOR2HS $T=739660 578040 0 180 $X=734080 $Y=572620
X3130 3003 2890 2977 2 1 XOR2HS $T=740280 547800 1 180 $X=734700 $Y=547420
X3131 2998 2977 3018 2 1 XOR2HS $T=737800 547800 1 0 $X=737800 $Y=542380
X3132 392 2921 3027 2 1 XOR2HS $T=739040 699000 0 0 $X=739040 $Y=698620
X3133 3008 2636 2999 2 1 XOR2HS $T=745240 618360 1 180 $X=739660 $Y=617980
X3134 2792 2799 3012 2 1 XOR2HS $T=739660 638520 1 0 $X=739660 $Y=633100
X3135 2906 2636 3019 2 1 XOR2HS $T=745860 578040 0 180 $X=740280 $Y=572620
X3136 2987 2792 3015 2 1 XOR2HS $T=740280 608280 1 0 $X=740280 $Y=602860
X3137 2697 3008 3042 2 1 XOR2HS $T=741520 628440 1 0 $X=741520 $Y=623020
X3138 2906 2624 3041 2 1 XOR2HS $T=749580 578040 1 180 $X=744000 $Y=577660
X3139 373 3031 3062 2 1 XOR2HS $T=744000 688920 1 0 $X=744000 $Y=683500
X3140 382 2921 3039 2 1 XOR2HS $T=744620 709080 1 0 $X=744620 $Y=703660
X3141 391 2921 3072 2 1 XOR2HS $T=745240 699000 0 0 $X=745240 $Y=698620
X3142 2906 2697 3078 2 1 XOR2HS $T=746480 578040 1 0 $X=746480 $Y=572620
X3143 367 376 3057 2 1 XOR2HS $T=747720 709080 0 0 $X=747720 $Y=708700
X3144 3068 382 417 2 1 XOR2HS $T=748960 719160 1 0 $X=748960 $Y=713740
X3145 2986 2715 3058 2 1 XOR2HS $T=750200 588120 1 0 $X=750200 $Y=582700
X3146 3074 2685 3102 2 1 XOR2HS $T=758260 638520 0 180 $X=752680 $Y=633100
X3147 392 418 3118 2 1 XOR2HS $T=753300 699000 1 0 $X=753300 $Y=693580
X3148 3074 2697 3120 2 1 XOR2HS $T=753920 618360 1 0 $X=753920 $Y=612940
X3149 376 418 3121 2 1 XOR2HS $T=753920 688920 1 0 $X=753920 $Y=683500
X3150 2649 2943 3126 2 1 XOR2HS $T=754540 588120 0 0 $X=754540 $Y=587740
X3151 2986 2697 3134 2 1 XOR2HS $T=755780 588120 1 0 $X=755780 $Y=582700
X3152 2943 2762 3135 2 1 XOR2HS $T=755780 598200 0 0 $X=755780 $Y=597820
X3153 2685 2943 3124 2 1 XOR2HS $T=755780 608280 1 0 $X=755780 $Y=602860
X3154 3074 2762 3136 2 1 XOR2HS $T=755780 628440 0 0 $X=755780 $Y=628060
X3155 2965 3123 3139 2 1 XOR2HS $T=756400 567960 1 0 $X=756400 $Y=562540
X3156 389 418 3137 2 1 XOR2HS $T=756400 688920 0 0 $X=756400 $Y=688540
X3157 3025 3054 3144 2 1 XOR2HS $T=757020 557880 0 0 $X=757020 $Y=557500
X3158 3128 3119 426 2 1 XOR2HS $T=759500 547800 1 0 $X=759500 $Y=542380
X3159 2822 2785 3164 2 1 XOR2HS $T=761360 628440 0 0 $X=761360 $Y=628060
X3160 2882 3142 3165 2 1 XOR2HS $T=761360 678840 0 0 $X=761360 $Y=678460
X3161 402 418 428 2 1 XOR2HS $T=761360 719160 1 0 $X=761360 $Y=713740
X3162 3005 2685 3171 2 1 XOR2HS $T=761980 608280 1 0 $X=761980 $Y=602860
X3163 400 418 3167 2 1 XOR2HS $T=761980 699000 0 0 $X=761980 $Y=698620
X3164 3068 400 3172 2 1 XOR2HS $T=761980 709080 1 0 $X=761980 $Y=703660
X3165 3068 402 3220 2 1 XOR2HS $T=768180 709080 0 0 $X=768180 $Y=708700
X3166 3173 3202 3242 2 1 XOR2HS $T=771900 688920 0 0 $X=771900 $Y=688540
X3167 3157 3016 3239 2 1 XOR2HS $T=772520 588120 0 0 $X=772520 $Y=587740
X3168 2750 3247 3262 2 1 XOR2HS $T=775000 658680 0 0 $X=775000 $Y=658300
X3169 3091 3266 3307 2 1 XOR2HS $T=781820 638520 1 0 $X=781820 $Y=633100
X3170 3204 3306 3340 2 1 XOR2HS $T=788020 628440 1 0 $X=788020 $Y=623020
X3171 3359 3357 438 2 1 XOR2HS $T=795460 547800 1 180 $X=789880 $Y=547420
X3172 3325 3310 3434 2 1 XOR2HS $T=801040 709080 0 0 $X=801040 $Y=708700
X3173 3460 3467 450 2 1 XOR2HS $T=811580 567960 0 180 $X=806000 $Y=562540
X3174 3440 3427 3470 2 1 XOR2HS $T=806620 638520 0 0 $X=806620 $Y=638140
X3175 3414 3434 3476 2 1 XOR2HS $T=807240 709080 0 0 $X=807240 $Y=708700
X3176 3471 3507 3518 2 1 XOR2HS $T=815920 648600 0 0 $X=815920 $Y=648220
X3177 3425 3513 460 2 1 XOR2HS $T=817780 588120 0 0 $X=817780 $Y=587740
X3178 458 459 3534 2 1 XOR2HS $T=819640 719160 1 0 $X=819640 $Y=713740
X3179 3289 3526 3540 2 1 XOR2HS $T=821500 648600 0 0 $X=821500 $Y=648220
X3180 3543 3550 3560 2 1 XOR2HS $T=826460 688920 1 0 $X=826460 $Y=683500
X3181 3472 3502 3563 2 1 XOR2HS $T=827080 678840 1 0 $X=827080 $Y=673420
X3182 3553 3548 3567 2 1 XOR2HS $T=828320 658680 0 0 $X=828320 $Y=658300
X3183 3595 3585 3573 2 1 XOR2HS $T=837620 678840 1 180 $X=832040 $Y=678460
X3184 3618 3613 3600 2 1 XOR2HS $T=842580 668760 1 180 $X=837000 $Y=668380
X3185 3612 3625 3657 2 1 XOR2HS $T=843820 608280 0 0 $X=843820 $Y=607900
X3186 3672 3661 3681 2 1 XOR2HS $T=848780 598200 0 0 $X=848780 $Y=597820
X3187 3673 3676 3683 2 1 XOR2HS $T=848780 688920 1 0 $X=848780 $Y=683500
X3188 3684 3685 3696 2 1 XOR2HS $T=852500 588120 1 0 $X=852500 $Y=582700
X3189 3634 3666 3698 2 1 XOR2HS $T=853740 598200 1 0 $X=853740 $Y=592780
X3190 3694 3692 500 2 1 XOR2HS $T=856220 547800 1 0 $X=856220 $Y=542380
X3191 3697 3688 3704 2 1 XOR2HS $T=856220 578040 1 0 $X=856220 $Y=572620
X3192 3652 498 501 2 1 XOR2HS $T=857460 557880 0 0 $X=857460 $Y=557500
X3193 3742 3735 3705 2 1 XOR2HS $T=869240 709080 0 180 $X=863660 $Y=703660
X3194 3761 3757 3737 2 1 XOR2HS $T=872340 628440 1 180 $X=866760 $Y=628060
X3195 3766 3752 3689 2 1 XOR2HS $T=872960 699000 0 180 $X=867380 $Y=693580
X3196 3876 3874 3840 2 1 XOR2HS $T=892180 699000 1 180 $X=886600 $Y=698620
X3197 535 3887 3876 2 1 XOR2HS $T=895280 709080 1 180 $X=889700 $Y=708700
X3198 3878 3888 3903 2 1 XOR2HS $T=891560 588120 1 0 $X=891560 $Y=582700
X3199 538 537 3887 2 1 XOR2HS $T=897140 719160 0 180 $X=891560 $Y=713740
X3200 3882 3902 3921 2 1 XOR2HS $T=894040 557880 0 0 $X=894040 $Y=557500
X3201 3957 3954 3810 2 1 XOR2HS $T=903340 678840 1 180 $X=897760 $Y=678460
X3202 534 541 3874 2 1 XOR2HS $T=899000 699000 0 0 $X=899000 $Y=698620
X3203 3966 3965 3928 2 1 XOR2HS $T=905200 567960 0 180 $X=899620 $Y=562540
X3204 3994 3978 4013 2 1 XOR2HS $T=908300 588120 1 0 $X=908300 $Y=582700
X3205 4027 4022 3930 2 1 XOR2HS $T=915120 628440 0 180 $X=909540 $Y=623020
X3206 4010 4004 4029 2 1 XOR2HS $T=910780 578040 0 0 $X=910780 $Y=577660
X3207 4014 3995 4039 2 1 XOR2HS $T=912640 598200 1 0 $X=912640 $Y=592780
X3208 4092 4033 4053 2 1 XOR2HS $T=924420 588120 0 180 $X=918840 $Y=582700
X3209 4096 4091 4060 2 1 XOR2HS $T=925040 578040 0 180 $X=919460 $Y=572620
X3210 4140 4142 580 2 1 XOR2HS $T=930000 547800 1 0 $X=930000 $Y=542380
X3211 4157 4158 4038 2 1 XOR2HS $T=934340 588120 1 0 $X=934340 $Y=582700
X3212 4195 4192 4179 2 1 XOR2HS $T=945500 688920 0 180 $X=939920 $Y=683500
X3213 4214 4209 4101 2 1 XOR2HS $T=950460 678840 0 180 $X=944880 $Y=673420
X3214 4257 4258 4268 2 1 XOR2HS $T=960380 678840 0 0 $X=960380 $Y=678460
X3215 867 876 1 842 887 828 2 MOAI1S $T=305040 658680 0 0 $X=305040 $Y=658300
X3216 997 1047 1 1024 1059 1091 2 MOAI1S $T=343480 648600 1 0 $X=343480 $Y=643180
X3217 1153 1257 1 1247 1231 1235 2 MOAI1S $T=373240 618360 0 180 $X=369520 $Y=612940
X3218 1257 1180 1 1274 1281 1271 2 MOAI1S $T=373860 618360 0 0 $X=373860 $Y=617980
X3219 1416 1344 1 1405 1344 1399 2 MOAI1S $T=402380 648600 0 180 $X=398660 $Y=643180
X3220 1153 1459 1 1443 1432 1410 2 MOAI1S $T=412300 618360 0 180 $X=408580 $Y=612940
X3221 1153 1408 1 1443 1483 1492 2 MOAI1S $T=413540 618360 1 0 $X=413540 $Y=612940
X3222 1488 88 1 1479 88 1463 2 MOAI1S $T=417260 709080 1 180 $X=413540 $Y=708700
X3223 1516 105 1 1531 1532 1539 2 MOAI1S $T=424700 699000 1 0 $X=424700 $Y=693580
X3224 2695 2703 1 2689 2718 2728 2 MOAI1S $T=697500 608280 1 0 $X=697500 $Y=602860
X3225 2677 2683 1 2737 2696 2720 2 MOAI1S $T=705560 608280 1 180 $X=701840 $Y=607900
X3226 2807 2779 1 2753 2721 2769 2 MOAI1S $T=712380 668760 1 180 $X=708660 $Y=668380
X3227 2781 2710 1 2773 2776 2729 2 MOAI1S $T=712380 688920 0 180 $X=708660 $Y=683500
X3228 2658 2841 1 2722 2826 2857 2 MOAI1S $T=722920 618360 1 180 $X=719200 $Y=617980
X3229 2852 2787 1 2735 2883 2865 2 MOAI1S $T=721060 578040 1 0 $X=721060 $Y=572620
X3230 2910 2799 1 2887 2859 2875 2 MOAI1S $T=726640 638520 0 180 $X=722920 $Y=633100
X3231 404 2968 1 2945 2949 2952 2 MOAI1S $T=735320 678840 1 180 $X=731600 $Y=678460
X3232 404 2991 1 2949 2995 3000 2 MOAI1S $T=742140 678840 1 180 $X=738420 $Y=678460
X3233 367 2994 1 409 410 3022 2 MOAI1S $T=741520 719160 1 0 $X=741520 $Y=713740
X3234 408 2994 1 410 3044 3048 2 MOAI1S $T=742760 709080 0 0 $X=742760 $Y=708700
X3235 3057 2994 1 410 3106 3122 2 MOAI1S $T=753300 709080 0 0 $X=753300 $Y=708700
X3236 3197 3191 1 3096 2701 3154 2 MOAI1S $T=770040 578040 1 180 $X=766320 $Y=577660
X3237 3191 3171 1 3170 2701 3212 2 MOAI1S $T=768180 598200 0 0 $X=768180 $Y=597820
X3238 2886 3191 1 3200 3177 3213 2 MOAI1S $T=768180 608280 0 0 $X=768180 $Y=607900
X3239 3134 3191 1 3200 3129 3244 2 MOAI1S $T=772520 578040 0 0 $X=772520 $Y=577660
X3240 3216 3191 1 3234 3200 3245 2 MOAI1S $T=772520 588120 1 0 $X=772520 $Y=582700
X3241 3132 3172 1 3237 3125 3263 2 MOAI1S $T=774380 709080 1 0 $X=774380 $Y=703660
X3242 3132 3220 1 3125 3206 3258 2 MOAI1S $T=775000 709080 0 0 $X=775000 $Y=708700
X3243 4335 4246 1 4335 4327 4325 2 MOAI1S $T=988280 608280 1 180 $X=984560 $Y=607900
X3244 4335 4198 1 4335 4319 4188 2 MOAI1S $T=988900 598200 1 180 $X=985180 $Y=597820
X3245 4335 4235 1 4335 4351 4349 2 MOAI1S $T=993240 618360 1 0 $X=993240 $Y=612940
X3246 628 4321 1 628 4370 4356 2 MOAI1S $T=993860 598200 0 0 $X=993860 $Y=597820
X3247 628 4353 1 628 4374 4373 2 MOAI1S $T=996340 598200 1 0 $X=996340 $Y=592780
X3248 680 688 681 2 1 ND2S $T=261640 608280 1 180 $X=259780 $Y=607900
X3249 691 713 683 2 1 ND2S $T=269700 618360 0 180 $X=267840 $Y=612940
X3250 708 726 710 2 1 ND2S $T=272180 578040 1 180 $X=270320 $Y=577660
X3251 779 838 824 2 1 ND2S $T=299460 608280 1 180 $X=297600 $Y=607900
X3252 869 905 893 2 1 ND2S $T=310620 648600 0 0 $X=310620 $Y=648220
X3253 851 935 927 2 1 ND2S $T=316820 638520 1 180 $X=314960 $Y=638140
X3254 22 947 18 2 1 ND2S $T=318680 547800 0 180 $X=316820 $Y=542380
X3255 951 957 915 2 1 ND2S $T=319920 557880 0 180 $X=318060 $Y=552460
X3256 922 1005 991 2 1 ND2S $T=325500 578040 0 0 $X=325500 $Y=577660
X3257 1026 1023 912 2 1 ND2S $T=334180 557880 0 180 $X=332320 $Y=552460
X3258 1119 1105 979 2 1 ND2S $T=349060 567960 1 180 $X=347200 $Y=567580
X3259 997 1095 1109 2 1 ND2S $T=347200 638520 0 0 $X=347200 $Y=638140
X3260 1210 1207 1031 2 1 ND2S $T=365800 557880 1 180 $X=363940 $Y=557500
X3261 1212 1270 1256 2 1 ND2S $T=371380 567960 0 0 $X=371380 $Y=567580
X3262 1256 1272 1172 2 1 ND2S $T=374480 567960 0 180 $X=372620 $Y=562540
X3263 1256 1285 1226 2 1 ND2S $T=376340 557880 1 180 $X=374480 $Y=557500
X3264 1181 1282 1260 2 1 ND2S $T=378200 688920 1 180 $X=376340 $Y=688540
X3265 1324 1349 1279 2 1 ND2S $T=388740 578040 0 180 $X=386880 $Y=572620
X3266 1352 1350 1310 2 1 ND2S $T=389980 547800 1 180 $X=388120 $Y=547420
X3267 1345 72 1325 2 1 ND2S $T=389360 547800 1 0 $X=389360 $Y=542380
X3268 1448 1416 1228 2 1 ND2S $T=408580 648600 1 0 $X=408580 $Y=643180
X3269 1295 1483 1408 2 1 ND2S $T=416640 618360 1 180 $X=414780 $Y=617980
X3270 84 1501 99 2 1 ND2S $T=415400 547800 0 0 $X=415400 $Y=547420
X3271 1542 1545 1541 2 1 ND2S $T=429040 638520 1 0 $X=429040 $Y=633100
X3272 1521 1569 1544 2 1 ND2S $T=431520 598200 0 0 $X=431520 $Y=597820
X3273 1648 1657 1639 2 1 ND2S $T=451360 628440 0 0 $X=451360 $Y=628060
X3274 136 1694 1707 2 1 ND2S $T=461900 719160 0 180 $X=460040 $Y=713740
X3275 1717 1711 1705 2 1 ND2S $T=465620 547800 1 180 $X=463760 $Y=547420
X3276 1694 1721 1747 2 1 ND2S $T=467480 709080 0 0 $X=467480 $Y=708700
X3277 1765 1763 1710 2 1 ND2S $T=473060 578040 0 180 $X=471200 $Y=572620
X3278 1799 1806 1748 2 1 ND2S $T=479880 578040 0 180 $X=478020 $Y=572620
X3279 1790 1796 1754 2 1 ND2S $T=479260 608280 1 0 $X=479260 $Y=602860
X3280 1812 1819 1766 2 1 ND2S $T=481740 588120 0 180 $X=479880 $Y=582700
X3281 1793 1820 1775 2 1 ND2S $T=480500 598200 1 0 $X=480500 $Y=592780
X3282 1840 1798 1718 2 1 ND2S $T=486080 557880 0 180 $X=484220 $Y=552460
X3283 2672 2650 2667 2 1 ND2S $T=689440 567960 1 0 $X=689440 $Y=562540
X3284 2733 2724 370 2 1 ND2S $T=701220 699000 0 0 $X=701220 $Y=698620
X3285 2671 2764 2761 2 1 ND2S $T=708660 588120 1 0 $X=708660 $Y=582700
X3286 2733 2759 374 2 1 ND2S $T=708660 719160 1 0 $X=708660 $Y=713740
X3287 2854 2889 2865 2 1 ND2S $T=724160 557880 1 180 $X=722300 $Y=557500
X3288 2854 2917 2871 2 1 ND2S $T=723540 557880 1 0 $X=723540 $Y=552460
X3289 2959 2963 2870 2 1 ND2S $T=732840 598200 1 0 $X=732840 $Y=592780
X3290 3012 3007 2910 2 1 ND2S $T=740280 628440 0 0 $X=740280 $Y=628060
X3291 3179 3189 3085 2 1 ND2S $T=766940 638520 0 180 $X=765080 $Y=633100
X3292 3181 3179 3005 2 1 ND2S $T=768800 608280 1 0 $X=768800 $Y=602860
X3293 3273 3265 3147 2 1 ND2S $T=780580 628440 1 180 $X=778720 $Y=628060
X3294 3367 3359 3360 2 1 ND2S $T=795460 557880 1 180 $X=793600 $Y=557500
X3295 3318 3387 3379 2 1 ND2S $T=798560 598200 0 180 $X=796700 $Y=592780
X3296 3390 3382 3397 2 1 ND2S $T=797940 578040 0 0 $X=797940 $Y=577660
X3297 3433 3421 3361 2 1 ND2S $T=804140 668760 0 180 $X=802280 $Y=663340
X3298 3408 3437 3430 2 1 ND2S $T=802900 678840 1 0 $X=802900 $Y=673420
X3299 3456 3495 3356 2 1 ND2S $T=814060 648600 0 0 $X=814060 $Y=648220
X3300 3464 3557 3551 2 1 ND2S $T=829560 699000 1 180 $X=827700 $Y=698620
X3301 3564 3584 3556 2 1 ND2S $T=833280 618360 0 0 $X=833280 $Y=617980
X3302 3593 3586 3582 2 1 ND2S $T=836380 688920 1 180 $X=834520 $Y=688540
X3303 3608 3595 3601 2 1 ND2S $T=836380 699000 1 0 $X=836380 $Y=693580
X3304 3614 3634 3602 2 1 ND2S $T=841340 588120 0 0 $X=841340 $Y=587740
X3305 3649 3618 3627 2 1 ND2S $T=845680 668760 1 180 $X=843820 $Y=668380
X3306 3665 3684 3669 2 1 ND2S $T=852500 578040 1 180 $X=850640 $Y=577660
X3307 3679 3673 3644 2 1 ND2S $T=850640 688920 0 0 $X=850640 $Y=688540
X3308 3691 3694 3674 2 1 ND2S $T=855600 547800 0 180 $X=853740 $Y=542380
X3309 3755 3728 3744 2 1 ND2S $T=866140 658680 1 0 $X=866140 $Y=653260
X3310 3736 3747 3745 2 1 ND2S $T=868620 547800 0 0 $X=868620 $Y=547420
X3311 3732 3761 3759 2 1 ND2S $T=869860 638520 1 0 $X=869860 $Y=633100
X3312 3777 3772 3743 2 1 ND2S $T=874200 557880 1 180 $X=872340 $Y=557500
X3313 3746 3780 3781 2 1 ND2S $T=876060 648600 1 0 $X=876060 $Y=643180
X3314 3795 3805 521 2 1 ND2S $T=880400 547800 1 180 $X=878540 $Y=547420
X3315 521 3812 3776 2 1 ND2S $T=881640 547800 0 180 $X=879780 $Y=542380
X3316 3845 3790 3826 2 1 ND2S $T=885360 658680 1 0 $X=885360 $Y=653260
X3317 3863 3856 3760 2 1 ND2S $T=889080 557880 0 180 $X=887220 $Y=552460
X3318 3875 3878 3854 2 1 ND2S $T=890940 588120 0 180 $X=889080 $Y=582700
X3319 3838 3860 3837 2 1 ND2S $T=891560 638520 0 180 $X=889700 $Y=633100
X3320 3883 3882 3815 2 1 ND2S $T=892180 567960 1 180 $X=890320 $Y=567580
X3321 3838 3900 3885 2 1 ND2S $T=891560 638520 0 0 $X=891560 $Y=638140
X3322 3894 3890 3841 2 1 ND2S $T=894040 557880 1 180 $X=892180 $Y=557500
X3323 3891 3899 3838 2 1 ND2S $T=894040 638520 0 180 $X=892180 $Y=633100
X3324 3896 3904 3889 2 1 ND2S $T=894660 598200 0 180 $X=892800 $Y=592780
X3325 3915 3869 3911 2 1 ND2S $T=894660 658680 0 0 $X=894660 $Y=658300
X3326 534 3933 541 2 1 ND2S $T=896520 699000 0 0 $X=896520 $Y=698620
X3327 3906 3916 3922 2 1 ND2S $T=897140 578040 1 0 $X=897140 $Y=572620
X3328 3922 3966 3822 2 1 ND2S $T=900860 578040 1 0 $X=900860 $Y=572620
X3329 3985 3994 3999 2 1 ND2S $T=907680 567960 0 0 $X=907680 $Y=567580
X3330 4002 3924 3982 2 1 ND2S $T=910160 648600 1 180 $X=908300 $Y=648220
X3331 3991 4014 4007 2 1 ND2S $T=910160 598200 1 0 $X=910160 $Y=592780
X3332 4034 3957 4026 2 1 ND2S $T=912640 678840 0 0 $X=912640 $Y=678460
X3333 4003 4010 4028 2 1 ND2S $T=913260 567960 1 0 $X=913260 $Y=562540
X3334 4009 4035 4019 2 1 ND2S $T=915120 638520 1 180 $X=913260 $Y=638140
X3335 4071 4027 4062 2 1 ND2S $T=918220 628440 0 0 $X=918220 $Y=628060
X3336 4070 4065 4094 2 1 ND2S $T=921940 678840 0 0 $X=921940 $Y=678460
X3337 4049 4096 4090 2 1 ND2S $T=923800 567960 1 0 $X=923800 $Y=562540
X3338 4097 4092 4108 2 1 ND2S $T=924420 588120 1 0 $X=924420 $Y=582700
X3339 4132 4104 4125 2 1 ND2S $T=926900 638520 1 0 $X=926900 $Y=633100
X3340 4135 4141 4150 2 1 ND2S $T=931240 628440 0 0 $X=931240 $Y=628060
X3341 4137 4140 4112 2 1 ND2S $T=931860 547800 0 0 $X=931860 $Y=547420
X3342 4153 4157 4117 2 1 ND2S $T=934340 588120 1 180 $X=932480 $Y=587740
X3343 4171 4176 4180 2 1 ND2S $T=939920 688920 1 180 $X=938060 $Y=688540
X3344 4187 4169 4184 2 1 ND2S $T=943020 638520 1 0 $X=943020 $Y=633100
X3345 4211 4195 4216 2 1 ND2S $T=948600 688920 1 0 $X=948600 $Y=683500
X3346 4229 4228 4224 2 1 ND2S $T=955420 557880 0 180 $X=953560 $Y=552460
X3347 4219 4242 4167 2 1 ND2S $T=956040 547800 1 180 $X=954180 $Y=547420
X3348 4250 4256 4259 2 1 ND2S $T=959140 709080 0 0 $X=959140 $Y=708700
X3349 4264 4274 609 2 1 ND2S $T=965960 688920 1 180 $X=964100 $Y=688540
X3350 4270 4271 4262 2 1 ND2S $T=965340 547800 0 0 $X=965340 $Y=547420
X3351 4305 4275 4283 2 1 ND2S $T=971540 547800 1 0 $X=971540 $Y=542380
X3352 4264 4334 4314 2 1 ND2S $T=981460 688920 1 180 $X=979600 $Y=688540
X3353 697 695 1 721 693 682 2 MOAI1H $T=265980 648600 1 0 $X=265980 $Y=643180
X3354 837 828 1 835 687 820 2 MOAI1H $T=302560 668760 0 180 $X=295120 $Y=663340
X3355 851 891 1 842 897 920 2 MOAI1H $T=307520 638520 1 0 $X=307520 $Y=633100
X3356 946 851 1 918 955 1002 2 MOAI1H $T=318060 628440 0 0 $X=318060 $Y=628060
X3357 962 868 1 866 949 984 2 MOAI1H $T=320540 658680 1 0 $X=320540 $Y=653260
X3358 1042 1000 1 1029 967 992 2 MOAI1H $T=337900 608280 0 180 $X=330460 $Y=602860
X3359 1266 1271 1 1265 1219 1255 2 MOAI1H $T=378820 608280 1 180 $X=371380 $Y=607900
X3360 1341 71 1 1359 1288 1376 2 MOAI1H $T=388740 699000 0 0 $X=388740 $Y=698620
X3361 2622 2684 1 2678 2702 2712 2 MOAI1H $T=692540 588120 0 0 $X=692540 $Y=587740
X3362 2777 2718 1 2798 2815 2718 2 MOAI1H $T=708660 608280 0 0 $X=708660 $Y=607900
X3363 2677 2811 1 2927 2934 2940 2 MOAI1H $T=724160 598200 1 0 $X=724160 $Y=592780
X3364 2999 2910 1 2970 3084 3056 2 MOAI1H $T=745240 618360 0 0 $X=745240 $Y=617980
X3365 698 685 1 2 INV2 $T=264740 588120 1 180 $X=262880 $Y=587740
X3366 696 708 1 2 INV2 $T=265980 598200 0 180 $X=264120 $Y=592780
X3367 750 734 1 2 INV2 $T=279000 608280 0 180 $X=277140 $Y=602860
X3368 707 752 1 2 INV2 $T=285820 588120 0 180 $X=283960 $Y=582700
X3369 779 783 1 2 INV2 $T=288920 608280 1 180 $X=287060 $Y=607900
X3370 931 893 1 2 INV2 $T=316200 648600 1 180 $X=314340 $Y=648220
X3371 998 995 1 2 INV2 $T=328600 688920 1 0 $X=328600 $Y=683500
X3372 1103 1024 1 2 INV2 $T=347820 648600 1 0 $X=347820 $Y=643180
X3373 1116 1065 1 2 INV2 $T=349060 638520 1 0 $X=349060 $Y=633100
X3374 1146 1103 1 2 INV2 $T=355260 638520 1 180 $X=353400 $Y=638140
X3375 1202 1116 1 2 INV2 $T=364560 638520 0 180 $X=362700 $Y=633100
X3376 1147 1234 1 2 INV2 $T=368900 638520 0 0 $X=368900 $Y=638140
X3377 950 1240 1 2 INV2 $T=369520 648600 0 0 $X=369520 $Y=648220
X3378 1362 1354 1 2 INV2 $T=391220 588120 0 180 $X=389360 $Y=582700
X3379 1348 1367 1 2 INV2 $T=393080 598200 1 0 $X=393080 $Y=592780
X3380 73 1322 1 2 INV2 $T=395560 709080 1 180 $X=393700 $Y=708700
X3381 1400 1017 1 2 INV2 $T=399280 608280 0 0 $X=399280 $Y=607900
X3382 1406 1236 1 2 INV2 $T=401140 618360 0 0 $X=401140 $Y=617980
X3383 74 82 1 2 INV2 $T=404240 557880 1 0 $X=404240 $Y=552460
X3384 91 1444 1 2 INV2 $T=411060 699000 1 180 $X=409200 $Y=698620
X3385 1475 1480 1 2 INV2 $T=414160 598200 1 0 $X=414160 $Y=592780
X3386 1513 1211 1 2 INV2 $T=424700 648600 1 0 $X=424700 $Y=643180
X3387 1558 1562 1 2 INV2 $T=432140 678840 0 0 $X=432140 $Y=678460
X3388 1614 1613 1 2 INV2 $T=442680 678840 1 180 $X=440820 $Y=678460
X3389 122 1637 1 2 INV2 $T=448880 709080 0 0 $X=448880 $Y=708700
X3390 160 1826 1 2 INV2 $T=486700 699000 0 0 $X=486700 $Y=698620
X3391 163 1838 1 2 INV2 $T=491660 699000 1 180 $X=489800 $Y=698620
X3392 168 1852 1 2 INV2 $T=494140 688920 0 0 $X=494140 $Y=688540
X3393 1971 1896 1 2 INV2 $T=518320 608280 0 0 $X=518320 $Y=607900
X3394 216 1984 1 2 INV2 $T=527000 547800 1 180 $X=525140 $Y=547420
X3395 2034 198 1 2 INV2 $T=530100 557880 1 0 $X=530100 $Y=552460
X3396 2021 2049 1 2 INV2 $T=532580 557880 1 0 $X=532580 $Y=552460
X3397 2034 2062 1 2 INV2 $T=535680 557880 1 0 $X=535680 $Y=552460
X3398 216 2085 1 2 INV2 $T=550560 547800 0 0 $X=550560 $Y=547420
X3399 216 237 1 2 INV2 $T=553040 547800 1 0 $X=553040 $Y=542380
X3400 2375 2273 1 2 INV2 $T=615040 608280 0 180 $X=613180 $Y=602860
X3401 2375 2406 1 2 INV2 $T=622480 578040 1 0 $X=622480 $Y=572620
X3402 2588 2613 1 2 INV2 $T=677040 608280 1 0 $X=677040 $Y=602860
X3403 2629 2673 1 2 INV2 $T=698740 598200 0 180 $X=696880 $Y=592780
X3404 2629 2714 1 2 INV2 $T=698740 598200 1 0 $X=698740 $Y=592780
X3405 2714 2663 1 2 INV2 $T=701220 598200 1 0 $X=701220 $Y=592780
X3406 2604 2713 1 2 INV2 $T=701840 618360 1 0 $X=701840 $Y=612940
X3407 2631 2758 1 2 INV2 $T=708040 628440 0 0 $X=708040 $Y=628060
X3408 2682 2799 1 2 INV2 $T=712380 638520 1 0 $X=712380 $Y=633100
X3409 2842 2680 1 2 INV2 $T=717960 578040 0 180 $X=716100 $Y=572620
X3410 2824 2838 1 2 INV2 $T=716720 688920 0 0 $X=716720 $Y=688540
X3411 381 2824 1 2 INV2 $T=717340 709080 1 0 $X=717340 $Y=703660
X3412 2853 2842 1 2 INV2 $T=719200 578040 0 0 $X=719200 $Y=577660
X3413 2722 2874 1 2 INV2 $T=720440 628440 0 0 $X=720440 $Y=628060
X3414 2874 2884 1 2 INV2 $T=722300 628440 0 0 $X=722300 $Y=628060
X3415 2874 2887 1 2 INV2 $T=724160 628440 0 0 $X=724160 $Y=628060
X3416 2683 2866 1 2 INV2 $T=726640 608280 0 180 $X=724780 $Y=602860
X3417 2837 2829 1 2 INV2 $T=728500 618360 0 180 $X=726640 $Y=612940
X3418 2910 2872 1 2 INV2 $T=726640 618360 0 0 $X=726640 $Y=617980
X3419 2929 2927 1 2 INV2 $T=728500 598200 0 0 $X=728500 $Y=597820
X3420 2929 2937 1 2 INV2 $T=728500 608280 1 0 $X=728500 $Y=602860
X3421 2671 2699 1 2 INV2 $T=729120 588120 1 0 $X=729120 $Y=582700
X3422 399 2949 1 2 INV2 $T=729740 709080 1 0 $X=729740 $Y=703660
X3423 2842 2953 1 2 INV2 $T=731600 578040 1 0 $X=731600 $Y=572620
X3424 2918 2960 1 2 INV2 $T=732840 608280 0 0 $X=732840 $Y=607900
X3425 2960 2959 1 2 INV2 $T=733460 598200 0 0 $X=733460 $Y=597820
X3426 2910 2912 1 2 INV2 $T=737800 628440 0 0 $X=737800 $Y=628060
X3427 412 3031 1 2 INV2 $T=749580 678840 0 0 $X=749580 $Y=678460
X3428 406 3125 1 2 INV2 $T=756400 719160 1 0 $X=756400 $Y=713740
X3429 2812 3202 1 2 INV2 $T=768800 699000 1 0 $X=768800 $Y=693580
X3430 2659 3200 1 2 INV2 $T=769420 588120 1 0 $X=769420 $Y=582700
X3431 3067 3235 1 2 INV2 $T=773140 598200 0 0 $X=773140 $Y=597820
X3432 3084 3271 1 2 INV2 $T=778100 608280 0 0 $X=778100 $Y=607900
X3433 3360 3386 1 2 INV2 $T=796080 557880 0 0 $X=796080 $Y=557500
X3434 3301 3395 1 2 INV2 $T=796700 648600 0 0 $X=796700 $Y=648220
X3435 3371 3403 1 2 INV2 $T=797940 658680 0 0 $X=797940 $Y=658300
X3436 3334 3433 1 2 INV2 $T=798560 668760 1 0 $X=798560 $Y=663340
X3437 3444 3441 1 2 INV2 $T=806000 678840 1 0 $X=806000 $Y=673420
X3438 3478 3455 1 2 INV2 $T=811580 628440 1 180 $X=809720 $Y=628060
X3439 3405 3465 1 2 INV2 $T=814060 678840 0 0 $X=814060 $Y=678460
X3440 3420 3492 1 2 INV2 $T=815300 618360 0 0 $X=815300 $Y=617980
X3441 3462 3506 1 2 INV2 $T=815920 608280 0 0 $X=815920 $Y=607900
X3442 3516 3493 1 2 INV2 $T=819020 628440 0 180 $X=817160 $Y=623020
X3443 3482 3527 1 2 INV2 $T=820260 668760 1 0 $X=820260 $Y=663340
X3444 166 3538 1 2 INV2 $T=824600 547800 0 0 $X=824600 $Y=547420
X3445 546 539 1 2 INV2 $T=902100 547800 0 180 $X=900240 $Y=542380
X3446 546 3951 1 2 INV2 $T=920080 547800 0 0 $X=920080 $Y=547420
X3447 574 4107 1 2 INV2 $T=926900 719160 0 180 $X=925040 $Y=713740
X3448 600 3718 1 2 INV2 $T=953560 638520 0 180 $X=951700 $Y=633100
X3449 611 4296 1 2 INV2 $T=970300 709080 1 180 $X=968440 $Y=708700
X3450 614 4301 1 2 INV2 $T=973400 719160 1 0 $X=973400 $Y=713740
X3451 4318 4314 1 2 INV2 $T=979600 699000 0 180 $X=977740 $Y=693580
X3452 4342 4329 1 2 INV2 $T=987660 709080 1 180 $X=985800 $Y=708700
X3453 4369 4340 1 2 INV2 $T=992000 688920 0 180 $X=990140 $Y=683500
X3454 4537 4523 1 2 INV2 $T=1074460 567960 1 0 $X=1074460 $Y=562540
X3455 1234 1173 1 2 BUF2 $T=372000 638520 0 180 $X=368900 $Y=633100
X3456 1071 1099 1 2 BUF2 $T=381300 688920 1 0 $X=381300 $Y=683500
X3457 1335 66 1 2 BUF2 $T=387500 719160 0 180 $X=384400 $Y=713740
X3458 1400 983 1 2 BUF2 $T=399900 618360 1 0 $X=399900 $Y=612940
X3459 1329 1433 1 2 BUF2 $T=407960 648600 0 0 $X=407960 $Y=648220
X3460 1536 1315 1 2 BUF2 $T=427800 628440 0 180 $X=424700 $Y=623020
X3461 1568 1422 1 2 BUF2 $T=442060 658680 1 180 $X=438960 $Y=658300
X3462 1590 124 1 2 BUF2 $T=447640 547800 1 180 $X=444540 $Y=547420
X3463 1635 1568 1 2 BUF2 $T=451360 658680 0 180 $X=448260 $Y=653260
X3464 1684 1525 1 2 BUF2 $T=457560 557880 0 180 $X=454460 $Y=552460
X3465 1699 1676 1 2 BUF2 $T=467480 648600 1 0 $X=467480 $Y=643180
X3466 1676 1851 1 2 BUF2 $T=484220 658680 1 0 $X=484220 $Y=653260
X3467 1854 1797 1 2 BUF2 $T=489180 648600 1 180 $X=486080 $Y=648220
X3468 1839 149 1 2 BUF2 $T=486080 709080 0 0 $X=486080 $Y=708700
X3469 1826 1858 1 2 BUF2 $T=486700 668760 0 0 $X=486700 $Y=668380
X3470 1863 1842 1 2 BUF2 $T=491040 628440 1 180 $X=487940 $Y=628060
X3471 1880 1839 1 2 BUF2 $T=499720 699000 0 180 $X=496620 $Y=693580
X3472 1902 1684 1 2 BUF2 $T=505300 557880 1 180 $X=502200 $Y=557500
X3473 1852 1895 1 2 BUF2 $T=504680 678840 1 0 $X=504680 $Y=673420
X3474 1938 1902 1 2 BUF2 $T=509020 567960 0 180 $X=505920 $Y=562540
X3475 1880 1940 1 2 BUF2 $T=508400 688920 0 0 $X=508400 $Y=688540
X3476 191 1938 1 2 BUF2 $T=512740 557880 0 0 $X=512740 $Y=557500
X3477 1851 2052 1 2 BUF2 $T=534440 658680 1 0 $X=534440 $Y=653260
X3478 1940 2039 1 2 BUF2 $T=535680 699000 0 0 $X=535680 $Y=698620
X3479 2062 247 1 2 BUF2 $T=552420 547800 0 0 $X=552420 $Y=547420
X3480 2046 2123 1 2 BUF2 $T=555520 578040 1 0 $X=555520 $Y=572620
X3481 2082 2375 1 2 BUF2 $T=615040 608280 1 0 $X=615040 $Y=602860
X3482 2338 2400 1 2 BUF2 $T=626820 567960 0 0 $X=626820 $Y=567580
X3483 2405 2526 1 2 BUF2 $T=651000 557880 0 0 $X=651000 $Y=557500
X3484 2557 2462 1 2 BUF2 $T=657820 668760 1 180 $X=654720 $Y=668380
X3485 2526 327 1 2 BUF2 $T=655340 557880 0 0 $X=655340 $Y=557500
X3486 2637 2626 1 2 BUF2 $T=683860 578040 1 180 $X=680760 $Y=577660
X3487 2663 2648 1 2 BUF2 $T=689440 608280 1 180 $X=686340 $Y=607900
X3488 2622 2671 1 2 BUF2 $T=689440 588120 0 0 $X=689440 $Y=587740
X3489 2618 2668 1 2 BUF2 $T=689440 638520 0 0 $X=689440 $Y=638140
X3490 2611 2618 1 2 BUF2 $T=693780 658680 1 180 $X=690680 $Y=658300
X3491 2641 2611 1 2 BUF2 $T=691300 678840 0 0 $X=691300 $Y=678460
X3492 357 2641 1 2 BUF2 $T=695640 709080 1 0 $X=695640 $Y=703660
X3493 2710 2733 1 2 BUF2 $T=706800 699000 0 180 $X=703700 $Y=693580
X3494 2627 2837 1 2 BUF2 $T=714860 608280 1 0 $X=714860 $Y=602860
X3495 2658 2910 1 2 BUF2 $T=723540 618360 0 0 $X=723540 $Y=617980
X3496 2884 2970 1 2 BUF2 $T=737180 618360 1 180 $X=734080 $Y=617980
X3497 2799 3008 1 2 BUF2 $T=740900 648600 1 0 $X=740900 $Y=643180
X3498 2987 3074 1 2 BUF2 $T=746480 608280 1 0 $X=746480 $Y=602860
X3499 3031 418 1 2 BUF2 $T=749580 688920 1 0 $X=749580 $Y=683500
X3500 3538 469 1 2 BUF2 $T=825220 557880 1 0 $X=825220 $Y=552460
X3501 3637 3547 1 2 BUF2 $T=843820 638520 1 180 $X=840720 $Y=638140
X3502 3547 3592 1 2 BUF2 $T=846920 638520 1 0 $X=846920 $Y=633100
X3503 3690 3637 1 2 BUF2 $T=854980 668760 1 0 $X=854980 $Y=663340
X3504 3592 3702 1 2 BUF2 $T=858700 618360 0 0 $X=858700 $Y=617980
X3505 3702 3783 1 2 BUF2 $T=870480 618360 1 0 $X=870480 $Y=612940
X3506 4202 589 1 2 BUF2 $T=953560 557880 1 180 $X=950460 $Y=557500
X3507 3718 4205 1 2 BUF2 $T=954180 588120 0 0 $X=954180 $Y=587740
X3508 4213 4041 1 2 BUF2 $T=964720 618360 0 180 $X=961620 $Y=612940
X3509 4213 4247 1 2 BUF2 $T=965340 618360 0 0 $X=965340 $Y=617980
X3510 4309 4213 1 2 BUF2 $T=975880 618360 1 180 $X=972780 $Y=617980
X3511 4255 4330 1 2 BUF2 $T=982080 567960 1 0 $X=982080 $Y=562540
X3512 4252 4255 1 2 BUF2 $T=983940 567960 0 0 $X=983940 $Y=567580
X3513 4313 4309 1 2 BUF2 $T=988280 628440 0 180 $X=985180 $Y=623020
X3514 4313 4367 1 2 BUF2 $T=990140 628440 1 0 $X=990140 $Y=623020
X3515 4330 619 1 2 BUF2 $T=993860 547800 0 180 $X=990760 $Y=542380
X3516 4345 4333 1 2 BUF2 $T=998820 658680 1 0 $X=998820 $Y=653260
X3517 4367 4345 1 2 BUF2 $T=1000680 638520 1 0 $X=1000680 $Y=633100
X3518 4359 637 1 2 BUF2 $T=1004400 547800 1 0 $X=1004400 $Y=542380
X3519 4428 4427 1 2 BUF2 $T=1026100 578040 0 0 $X=1026100 $Y=577660
X3520 4490 4438 1 2 BUF2 $T=1048420 598200 1 180 $X=1045320 $Y=597820
X3521 4475 4452 1 2 BUF2 $T=1052760 709080 0 180 $X=1049660 $Y=703660
X3522 4452 4487 1 2 BUF2 $T=1050280 688920 1 0 $X=1050280 $Y=683500
X3523 653 4475 1 2 BUF2 $T=1054620 709080 1 180 $X=1051520 $Y=708700
X3524 4510 4490 1 2 BUF2 $T=1057100 588120 0 180 $X=1054000 $Y=582700
X3525 4487 4514 1 2 BUF2 $T=1063920 678840 0 180 $X=1060820 $Y=673420
X3526 4517 4566 1 2 BUF2 $T=1078180 688920 0 0 $X=1078180 $Y=688540
X3527 4514 4562 1 2 BUF2 $T=1081900 668760 0 0 $X=1081900 $Y=668380
X3528 4569 4601 1 2 BUF2 $T=1089960 567960 1 0 $X=1089960 $Y=562540
X3529 4601 4604 1 2 BUF2 $T=1098640 567960 1 0 $X=1098640 $Y=562540
X3530 4618 4600 1 2 BUF2 $T=1106700 638520 0 180 $X=1103600 $Y=633100
X3531 4604 4613 1 2 BUF2 $T=1107940 588120 0 180 $X=1104840 $Y=582700
X3532 4600 4594 1 2 BUF2 $T=1106080 648600 1 0 $X=1106080 $Y=643180
X3533 4591 4618 1 2 BUF2 $T=1114140 628440 1 0 $X=1114140 $Y=623020
X3534 1516 81 106 2 107 110 1 AO22 $T=424080 719160 1 0 $X=424080 $Y=713740
X3535 686 680 1 2 INV3 $T=259780 618360 0 180 $X=257300 $Y=612940
X3536 931 866 1 2 INV3 $T=326120 648600 0 0 $X=326120 $Y=648220
X3537 1103 1016 1 2 INV3 $T=347820 658680 0 180 $X=345340 $Y=653260
X3538 1165 931 1 2 INV3 $T=358360 648600 0 180 $X=355880 $Y=643180
X3539 1306 786 1 2 INV3 $T=381300 658680 1 0 $X=381300 $Y=653260
X3540 189 1952 1 2 INV3 $T=511500 588120 0 0 $X=511500 $Y=587740
X3541 1963 2034 1 2 INV3 $T=537540 567960 1 180 $X=535060 $Y=567580
X3542 2082 2096 1 2 INV3 $T=541880 598200 0 0 $X=541880 $Y=597820
X3543 291 2402 1 2 INV3 $T=615040 688920 1 0 $X=615040 $Y=683500
X3544 292 2082 1 2 INV3 $T=615040 688920 0 0 $X=615040 $Y=688540
X3545 2633 2629 1 2 INV3 $T=683240 588120 1 180 $X=680760 $Y=587740
X3546 2659 2678 1 2 INV3 $T=698120 588120 1 0 $X=698120 $Y=582700
X3547 2815 2918 1 2 INV3 $T=732840 608280 1 180 $X=730360 $Y=607900
X3548 3473 3436 1 2 INV3 $T=810340 578040 0 0 $X=810340 $Y=577660
X3549 600 4418 1 2 INV3 $T=1011220 658680 0 180 $X=1008740 $Y=653260
X3550 4484 4537 1 2 INV3 $T=1058960 567960 0 0 $X=1058960 $Y=567580
X3551 4537 4569 1 2 INV3 $T=1078180 567960 1 0 $X=1078180 $Y=562540
X3552 4570 4591 1 2 INV3 $T=1086240 628440 1 0 $X=1086240 $Y=623020
X3553 1153 867 1 2 BUF6 $T=357120 618360 0 180 $X=349680 $Y=612940
X3554 1453 1306 1 2 BUF6 $T=411060 658680 0 180 $X=403620 $Y=653260
X3555 1378 1344 1 2 BUF6 $T=417260 628440 1 0 $X=417260 $Y=623020
X3556 1637 86 1 2 BUF6 $T=448880 709080 1 180 $X=441440 $Y=708700
X3557 1691 1635 1 2 BUF6 $T=465000 668760 0 0 $X=465000 $Y=668380
X3558 1764 1691 1 2 BUF6 $T=474300 688920 0 180 $X=466860 $Y=683500
X3559 1927 1955 1 2 BUF6 $T=522660 588120 1 0 $X=522660 $Y=582700
X3560 1952 2046 1 2 BUF6 $T=537540 567960 0 0 $X=537540 $Y=567580
X3561 2049 244 1 2 BUF6 $T=544980 557880 1 0 $X=544980 $Y=552460
X3562 2322 2057 1 2 BUF6 $T=608220 598200 0 0 $X=608220 $Y=597820
X3563 2391 2322 1 2 BUF6 $T=629300 618360 1 180 $X=621860 $Y=617980
X3564 2733 369 1 2 BUF6 $T=708660 719160 0 180 $X=701220 $Y=713740
X3565 3356 3351 1 2 BUF6 $T=819640 678840 1 0 $X=819640 $Y=673420
X3566 4418 4437 1 2 BUF6 $T=1023620 648600 1 0 $X=1023620 $Y=643180
X3567 4437 4474 1 2 BUF6 $T=1037260 628440 0 0 $X=1037260 $Y=628060
X3568 4427 4484 1 2 BUF6 $T=1042840 578040 1 0 $X=1042840 $Y=572620
X3569 4474 4508 1 2 BUF6 $T=1054620 638520 0 180 $X=1047180 $Y=633100
X3570 4508 4534 1 2 BUF6 $T=1063920 628440 0 0 $X=1063920 $Y=628060
X3571 864 1 869 866 837 861 2 OAI22S $T=306280 668760 1 180 $X=302560 $Y=668380
X3572 861 1 869 866 877 881 2 OAI22S $T=303180 678840 1 0 $X=303180 $Y=673420
X3573 1051 1 1020 1024 1019 1011 2 OAI22S $T=336040 638520 0 180 $X=332320 $Y=633100
X3574 1011 1 1020 1024 936 1021 2 OAI22S $T=332320 638520 0 0 $X=332320 $Y=638140
X3575 1065 1 1021 1024 878 1037 2 OAI22S $T=338520 648600 0 180 $X=334800 $Y=643180
X3576 1059 1 1020 1024 1054 1051 2 OAI22S $T=340380 638520 0 180 $X=336660 $Y=633100
X3577 1086 1 1065 1016 1098 1104 2 OAI22S $T=344100 668760 0 0 $X=344100 $Y=668380
X3578 1050 1 1065 1016 964 1076 2 OAI22S $T=347820 678840 1 180 $X=344100 $Y=678460
X3579 1104 1 1065 1146 1139 1164 2 OAI22S $T=354020 638520 1 0 $X=354020 $Y=633100
X3580 1164 1 1202 1146 1227 1248 2 OAI22S $T=366420 628440 0 0 $X=366420 $Y=628060
X3581 1221 1 1240 1252 1253 1165 2 OAI22S $T=368900 648600 1 0 $X=368900 $Y=643180
X3582 1202 1 1248 1146 1259 1258 2 OAI22S $T=375720 628440 1 180 $X=372000 $Y=628060
X3583 69 1 70 66 1341 75 2 OAI22S $T=388120 719160 1 0 $X=388120 $Y=713740
X3584 1473 1 1240 1389 1518 1530 2 OAI22S $T=422220 628440 0 0 $X=422220 $Y=628060
X3585 1394 1 121 1335 1617 128 2 OAI22S $T=444540 719160 1 0 $X=444540 $Y=713740
X3586 2712 1 2699 2678 2744 2748 2 OAI22S $T=701220 588120 1 0 $X=701220 $Y=582700
X3587 2793 1 2800 2776 2807 2831 2 OAI22S $T=711760 678840 1 0 $X=711760 $Y=673420
X3588 2773 1 2800 2776 2763 2793 2 OAI22S $T=711760 678840 0 0 $X=711760 $Y=678460
X3589 2813 1 379 381 2840 385 2 OAI22S $T=714860 709080 0 0 $X=714860 $Y=708700
X3590 2803 1 2701 2843 2849 2699 2 OAI22S $T=716100 588120 1 0 $X=716100 $Y=582700
X3591 2831 1 2800 2776 2836 2880 2 OAI22S $T=716720 678840 1 0 $X=716720 $Y=673420
X3592 2880 1 2800 2838 2903 2907 2 OAI22S $T=722300 678840 1 0 $X=722300 $Y=673420
X3593 2914 1 2800 2838 2904 2885 2 OAI22S $T=727880 688920 1 180 $X=724160 $Y=688540
X3594 2859 1 2912 2887 2896 2947 2 OAI22S $T=725400 638520 0 0 $X=725400 $Y=638140
X3595 2815 1 2955 2829 2923 2937 2 OAI22S $T=734080 618360 0 180 $X=730360 $Y=612940
X3596 2947 1 2912 2887 2938 2972 2 OAI22S $T=730980 638520 0 0 $X=730980 $Y=638140
X3597 2984 1 2699 2678 2966 2843 2 OAI22S $T=736560 588120 0 180 $X=732840 $Y=582700
X3598 2872 1 2983 2884 2975 2848 2 OAI22S $T=737800 628440 0 180 $X=734080 $Y=623020
X3599 2872 1 2989 2970 2993 3004 2 OAI22S $T=735940 618360 1 0 $X=735940 $Y=612940
X3600 2972 1 2912 2887 3030 3038 2 OAI22S $T=740900 638520 0 0 $X=740900 $Y=638140
X3601 2912 1 3056 3046 3067 2970 2 OAI22S $T=745860 628440 0 0 $X=745860 $Y=628060
X3602 2912 1 3038 3070 3076 2970 2 OAI22S $T=747100 638520 1 0 $X=747100 $Y=633100
X3603 2815 1 3083 2937 3107 3109 2 OAI22S $T=752060 608280 0 0 $X=752060 $Y=607900
X3604 3125 1 3141 424 3138 3106 2 OAI22S $T=762600 709080 1 180 $X=758880 $Y=708700
X3605 3162 1 3096 3151 3148 2701 2 OAI22S $T=765080 578040 1 180 $X=761360 $Y=577660
X3606 3170 1 3162 3200 3224 3193 2 OAI22S $T=770040 598200 1 0 $X=770040 $Y=592780
X3607 816 2 766 803 5 1 10 FA1S $T=290780 547800 1 0 $X=290780 $Y=542380
X3608 8 2 749 12 6 1 889 FA1S $T=295120 547800 0 0 $X=295120 $Y=547420
X3609 865 2 833 815 9 1 913 FA1S $T=299460 557880 1 0 $X=299460 $Y=552460
X3610 884 2 754 853 13 1 940 FA1S $T=302560 557880 0 0 $X=302560 $Y=557500
X3611 909 2 857 908 17 1 943 FA1S $T=306900 567960 1 0 $X=306900 $Y=562540
X3612 973 2 917 953 27 1 1008 FA1S $T=318680 557880 0 0 $X=318680 $Y=557500
X3613 1040 2 1052 982 35 1 990 FA1S $T=340380 547800 1 180 $X=328600 $Y=547420
X3614 1041 2 1009 1006 36 1 1032 FA1S $T=331080 567960 1 0 $X=331080 $Y=562540
X3615 1074 2 1096 1043 41 1 1113 FA1S $T=337900 557880 0 0 $X=337900 $Y=557500
X3616 1134 2 1123 1110 49 1 1170 FA1S $T=348440 547800 1 0 $X=348440 $Y=542380
X3617 1218 2 1192 1196 56 1 1262 FA1S $T=362080 547800 0 0 $X=362080 $Y=547420
X3618 1316 2 1370 1333 68 1 1374 FA1S $T=385020 557880 1 0 $X=385020 $Y=552460
X3619 1360 2 1392 1401 90 1 1450 FA1S $T=398040 547800 0 0 $X=398040 $Y=547420
X3620 1669 2 1551 1616 135 1 1706 FA1S $T=451360 557880 0 0 $X=451360 $Y=557500
X3621 1697 2 1714 1672 133 1 1733 FA1S $T=456320 598200 1 0 $X=456320 $Y=592780
X3622 1701 2 1673 1724 139 1 1735 FA1S $T=456940 578040 0 0 $X=456940 $Y=577660
X3623 1702 2 1698 1677 134 1 1760 FA1S $T=456940 598200 0 0 $X=456940 $Y=597820
X3624 1712 2 1692 1722 144 1 1685 FA1S $T=469340 588120 1 180 $X=457560 $Y=587740
X3625 1708 2 1696 1732 146 1 1695 FA1S $T=472440 567960 1 180 $X=460660 $Y=567580
X3626 2816 2 2791 2795 2896 1 2897 FA1S $T=709900 648600 1 0 $X=709900 $Y=643180
X3627 3594 2 481 3570 2377 1 3640 FA1S $T=832040 578040 1 0 $X=832040 $Y=572620
X3628 3599 2 484 468 475 1 3604 FA1S $T=833280 719160 1 0 $X=833280 $Y=713740
X3629 480 2 477 3580 3531 1 486 FA1S $T=834520 547800 1 0 $X=834520 $Y=542380
X3630 3655 2 3656 487 491 1 3623 FA1S $T=854980 709080 1 180 $X=843200 $Y=708700
X3631 3708 2 3725 497 3709 1 3671 FA1S $T=866140 699000 1 180 $X=854360 $Y=698620
X3632 3710 2 499 3706 3616 1 513 FA1S $T=858080 557880 1 0 $X=858080 $Y=552460
X3633 3720 2 503 3707 3588 1 3739 FA1S $T=860560 567960 0 0 $X=860560 $Y=567580
X3634 3740 2 507 3726 3561 1 3779 FA1S $T=863660 578040 1 0 $X=863660 $Y=572620
X3635 3753 2 517 3778 3611 1 3765 FA1S $T=865520 588120 0 0 $X=865520 $Y=587740
X3636 3774 2 3748 519 3734 1 3729 FA1S $T=877920 668760 1 180 $X=866140 $Y=668380
X3637 3799 2 3764 526 3758 1 3763 FA1S $T=882880 688920 1 180 $X=871100 $Y=688540
X3638 3831 2 527 3859 3568 1 3855 FA1S $T=878540 598200 0 0 $X=878540 $Y=597820
X3639 3839 2 3870 531 3802 1 3814 FA1S $T=892180 668760 1 180 $X=880400 $Y=668380
X3640 3865 2 3919 540 3727 1 3850 FA1S $T=898380 668760 0 180 $X=886600 $Y=663340
X3641 3923 2 532 3961 3792 1 3979 FA1S $T=893420 598200 0 0 $X=893420 $Y=597820
X3642 3934 2 4056 548 3722 1 3872 FA1S $T=905200 678840 0 180 $X=893420 $Y=673420
X3643 3953 2 4020 558 3719 1 3937 FA1S $T=912020 668760 1 180 $X=900240 $Y=668380
X3644 3992 2 550 4021 3615 1 4017 FA1S $T=903960 557880 1 0 $X=903960 $Y=552460
X3645 4011 2 4006 565 3682 1 3968 FA1S $T=918220 658680 1 180 $X=906440 $Y=658300
X3646 557 2 561 3986 3578 1 4025 FA1S $T=907060 547800 0 0 $X=907060 $Y=547420
X3647 4057 2 4133 572 3716 1 4037 FA1S $T=927520 658680 0 180 $X=915740 $Y=653260
X3648 4128 2 4178 584 3662 1 4000 FA1S $T=935580 658680 1 180 $X=923800 $Y=658300
X3649 4145 2 4170 588 3713 1 4110 FA1S $T=939300 648600 1 180 $X=927520 $Y=648220
X3650 4166 2 4221 593 3703 1 4151 FA1S $T=946120 658680 0 180 $X=934340 $Y=653260
X3651 4084 2 4231 603 3641 1 4191 FA1S $T=954800 648600 1 180 $X=943020 $Y=648220
X3652 4199 2 4230 599 3701 1 4175 FA1S $T=955420 648600 0 180 $X=943640 $Y=643180
X3653 4336 2 4327 4246 4358 1 4635 FA1S $T=981460 618360 1 0 $X=981460 $Y=612940
X3654 4358 2 4351 4235 4377 1 4636 FA1S $T=991380 608280 0 0 $X=991380 $Y=607900
X3655 4377 2 4370 4321 4383 1 4637 FA1S $T=995720 608280 1 0 $X=995720 $Y=602860
X3656 4383 2 4374 4353 635 1 4638 FA1S $T=998200 598200 0 0 $X=998200 $Y=597820
X3657 1299 1153 1 2 INV4 $T=380060 618360 0 180 $X=376960 $Y=612940
X3658 1971 1863 1 2 INV4 $T=516460 618360 0 180 $X=513360 $Y=612940
X3659 2021 1989 1 2 INV4 $T=527000 547800 0 0 $X=527000 $Y=547420
X3660 1988 2021 1 2 INV4 $T=532580 557880 1 180 $X=529480 $Y=557500
X3661 295 2410 1 2 INV4 $T=618760 688920 0 0 $X=618760 $Y=688540
X3662 600 638 1 2 INV4 $T=1009980 598200 0 0 $X=1009980 $Y=597820
X3663 4570 4551 1 2 INV4 $T=1082520 618360 0 180 $X=1079420 $Y=612940
X3664 4534 4570 1 2 INV4 $T=1083140 628440 0 180 $X=1080040 $Y=623020
X3665 767 772 1 768 2 OR2T $T=289540 598200 0 180 $X=283340 $Y=592780
X3666 813 840 1 750 2 OR2T $T=300700 598200 1 180 $X=294500 $Y=597820
X3667 1347 1287 1 1324 2 OR2T $T=388740 588120 1 180 $X=382540 $Y=587740
X3668 1353 976 1 1326 2 OR2T $T=391220 618360 0 180 $X=385020 $Y=612940
X3669 1409 1418 1 1426 2 OR2T $T=399900 688920 1 0 $X=399900 $Y=683500
X3670 1444 83 1 1376 2 OR2T $T=409200 699000 1 180 $X=403000 $Y=698620
X3671 98 1468 1 102 2 OR2T $T=417880 719160 1 0 $X=417880 $Y=713740
X3672 1579 1526 1 1600 2 OR2T $T=435240 618360 0 0 $X=435240 $Y=617980
X3673 4227 4251 1 4238 2 OR2T $T=957280 699000 0 0 $X=957280 $Y=698620
X3674 1236 1281 1365 1201 2 1378 1 AOI13HS $T=392460 628440 1 0 $X=392460 $Y=623020
X3675 2713 2737 2745 2628 2 2718 1 AOI13HS $T=703700 618360 1 0 $X=703700 $Y=612940
X3676 3657 2 3680 3681 3699 1 NR3 $T=850020 608280 1 0 $X=850020 $Y=602860
X3677 45 952 1081 1 2 47 OA12 $T=344720 547800 1 0 $X=344720 $Y=542380
X3678 1294 1146 1283 1 2 1321 OA12 $T=378200 628440 0 0 $X=378200 $Y=628060
X3679 1540 1389 1545 1 2 1550 OA12 $T=427180 628440 0 0 $X=427180 $Y=628060
X3680 1563 1581 1544 1 2 1573 OA12 $T=438340 608280 0 180 $X=434620 $Y=602860
X3681 1636 1614 1632 1 2 1623 OA12 $T=448260 678840 1 180 $X=444540 $Y=678460
X3682 1642 1627 1639 1 2 1610 OA12 $T=450120 628440 0 180 $X=446400 $Y=623020
X3683 1637 1335 1650 1 2 1664 OA12 $T=448880 709080 1 0 $X=448880 $Y=703660
X3684 130 1335 132 1 2 1667 OA12 $T=451980 719160 1 0 $X=451980 $Y=713740
X3685 1719 141 1694 1 2 1690 OA12 $T=466240 709080 1 180 $X=462520 $Y=708700
X3686 2655 2670 2667 1 2 361 OA12 $T=690060 557880 0 0 $X=690060 $Y=557500
X3687 2701 2760 2764 1 2 2717 OA12 $T=709900 578040 1 180 $X=706180 $Y=577660
X3688 2983 2970 3007 1 2 3016 OA12 $T=737800 628440 1 0 $X=737800 $Y=623020
X3689 3152 3158 3186 1 2 3229 OA12 $T=770040 658680 1 0 $X=770040 $Y=653260
X3690 3230 3200 3240 1 2 3251 OA12 $T=773760 608280 0 0 $X=773760 $Y=607900
X3691 3469 3418 3400 1 2 3494 OA12 $T=810340 638520 1 0 $X=810340 $Y=633100
X3692 3468 3448 3438 1 2 3496 OA12 $T=810340 688920 1 0 $X=810340 $Y=683500
X3693 4035 4022 4032 1 2 3996 OA12 $T=916980 638520 0 180 $X=913260 $Y=633100
X3694 869 984 1 866 1117 1124 2 OAI22H $T=344100 648600 0 0 $X=344100 $Y=648220
X3695 2800 2851 1 2838 2839 2780 2 OAI22H $T=722920 688920 0 180 $X=715480 $Y=683500
X3696 2872 2749 1 2722 2844 2809 2 OAI22H $T=723540 628440 0 180 $X=716100 $Y=623020
X3697 1383 3 1415 1121 1 2 QDFFRBP $T=410440 588120 0 180 $X=398040 $Y=582700
X3698 1425 3 1415 1371 1 2 QDFFRBP $T=411060 588120 1 180 $X=398660 $Y=587740
X3699 1455 3 1415 1400 1 2 QDFFRBP $T=411060 598200 1 180 $X=398660 $Y=597820
X3700 1529 11 1422 89 1 2 QDFFRBP $T=422840 668760 0 180 $X=410440 $Y=663340
X3701 1491 11 1422 112 1 2 QDFFRBP $T=420980 668760 0 0 $X=420980 $Y=668380
X3702 1586 116 1481 1378 1 2 QDFFRBP $T=440200 588120 1 180 $X=427800 $Y=587740
X3703 1554 11 1568 111 1 2 QDFFRBP $T=442060 668760 0 180 $X=429660 $Y=663340
X3704 1597 116 1641 1566 1 2 QDFFRBP $T=442680 588120 0 0 $X=442680 $Y=587740
X3705 1689 11 1635 108 1 2 QDFFRBP $T=463140 668760 1 180 $X=450740 $Y=668380
X3706 1740 11 1699 1223 1 2 QDFFRBP $T=469340 638520 0 180 $X=456940 $Y=633100
X3707 1741 11 1757 145 1 2 QDFFRBP $T=480500 699000 1 180 $X=468100 $Y=698620
X3708 2554 2290 2613 2627 1 2 QDFFRBP $T=668980 598200 0 0 $X=668980 $Y=597820
X3709 2599 2290 2589 2631 1 2 QDFFRBP $T=671460 618360 1 0 $X=671460 $Y=612940
X3710 2566 250 2613 2637 1 2 QDFFRBP $T=672080 578040 1 0 $X=672080 $Y=572620
X3711 2602 250 2613 2633 1 2 QDFFRBP $T=672080 588120 1 0 $X=672080 $Y=582700
X3712 2646 271 2641 2710 1 2 QDFFRBP $T=686340 688920 1 0 $X=686340 $Y=683500
X3713 2660 271 2641 365 1 2 QDFFRBP $T=688820 699000 0 0 $X=688820 $Y=698620
X3714 2661 271 357 367 1 2 QDFFRBP $T=688820 709080 0 0 $X=688820 $Y=708700
X3715 360 271 357 366 1 2 QDFFRBP $T=688820 719160 1 0 $X=688820 $Y=713740
X3716 740 3 738 2 1 833 QDFFRBS $T=285200 557880 0 0 $X=285200 $Y=557500
X3717 761 3 738 2 1 857 QDFFRBS $T=290780 567960 1 0 $X=290780 $Y=562540
X3718 1723 11 1676 2 1 1155 QDFFRBS $T=465000 648600 0 180 $X=453220 $Y=643180
X3719 4101 4080 4047 2 1 4006 QDFFRBS $T=925660 668760 0 180 $X=913880 $Y=663340
X3720 4179 4080 4047 2 1 4020 QDFFRBS $T=942400 668760 1 180 $X=930620 $Y=668380
X3721 4306 4080 4239 2 1 4231 QDFFRBS $T=980220 668760 0 180 $X=968440 $Y=663340
X3722 1826 155 1 154 1838 2 1778 1343 1852 OAI222S $T=482360 678840 0 0 $X=482360 $Y=678460
X3723 1826 158 1 159 1838 2 156 1411 1852 OAI222S $T=484220 688920 0 0 $X=484220 $Y=688540
X3724 1858 162 1 1879 1883 2 1856 1674 1895 OAI222S $T=492280 668760 1 0 $X=492280 $Y=663340
X3725 1865 1843 1 1847 1878 2 1864 1740 1894 OAI222S $T=495380 638520 1 0 $X=495380 $Y=633100
X3726 1826 176 1 1898 1838 2 1889 1338 1852 OAI222S $T=502200 678840 0 180 $X=496620 $Y=673420
X3727 1858 1901 1 1868 1883 2 1876 1628 1895 OAI222S $T=498480 648600 1 0 $X=498480 $Y=643180
X3728 1906 1927 1 1853 1931 2 1910 182 1942 OAI222S $T=504680 588120 0 0 $X=504680 $Y=587740
X3729 1922 1927 1 1903 1931 2 1939 188 1942 OAI222S $T=506540 598200 1 0 $X=506540 $Y=592780
X3730 1865 1928 1 1908 1878 2 1918 1809 1894 OAI222S $T=506540 638520 1 0 $X=506540 $Y=633100
X3731 1858 1937 1 1945 1883 2 1950 1407 1895 OAI222S $T=509020 668760 0 0 $X=509020 $Y=668380
X3732 1865 1960 1 1926 1878 2 1935 1816 1894 OAI222S $T=517080 638520 1 180 $X=511500 $Y=638140
X3733 1949 1955 1 1915 1963 2 1966 193 1988 OAI222S $T=512120 588120 1 0 $X=512120 $Y=582700
X3734 1943 198 1 1984 1987 2 1992 199 1989 OAI222S $T=516460 557880 1 0 $X=516460 $Y=552460
X3735 1858 202 1 1990 1883 2 1979 1668 1895 OAI222S $T=522040 668760 1 180 $X=516460 $Y=668380
X3736 1958 1955 1 1823 1963 2 1985 206 1988 OAI222S $T=517080 588120 0 0 $X=517080 $Y=587740
X3737 1865 1982 1 1961 1878 2 1997 1808 1894 OAI222S $T=517080 638520 0 0 $X=517080 $Y=638140
X3738 207 1984 1 187 198 2 1978 205 1989 OAI222S $T=525140 547800 1 180 $X=519560 $Y=547420
X3739 1858 2000 1 1998 1883 2 2010 1454 1895 OAI222S $T=520800 658680 0 0 $X=520800 $Y=658300
X3740 2003 1984 1 174 198 2 2019 209 1989 OAI222S $T=523280 557880 1 0 $X=523280 $Y=552460
X3741 1927 1910 1 1906 1931 2 2033 215 1942 OAI222S $T=526380 598200 1 0 $X=526380 $Y=592780
X3742 2032 1955 1 1835 1963 2 2036 218 1988 OAI222S $T=527620 588120 0 0 $X=527620 $Y=587740
X3743 1955 1992 1 1987 1963 2 2043 221 1988 OAI222S $T=529480 567960 0 0 $X=529480 $Y=567580
X3744 1955 1966 1 1949 1963 2 2050 225 1988 OAI222S $T=531340 588120 1 0 $X=531340 $Y=582700
X3745 1927 1939 1 1922 1931 2 2080 232 1942 OAI222S $T=537540 598200 1 0 $X=537540 $Y=592780
X3746 1984 1978 1 207 2062 2 2084 229 2049 OAI222S $T=538780 557880 1 0 $X=538780 $Y=552460
X3747 213 2062 1 2049 2094 2 222 236 2085 OAI222S $T=548080 557880 1 180 $X=542500 $Y=557500
X3748 1927 1985 1 1958 2096 2 2095 242 1942 OAI222S $T=543740 588120 0 0 $X=543740 $Y=587740
X3749 2110 2036 1 2032 2096 2 2116 246 2057 OAI222S $T=547460 598200 1 0 $X=547460 $Y=592780
X3750 2085 2019 1 2003 247 2 2128 248 244 OAI222S $T=552420 557880 1 0 $X=552420 $Y=552460
X3751 2085 231 1 203 247 2 2133 253 244 OAI222S $T=553660 557880 0 0 $X=553660 $Y=557500
X3752 2110 2219 1 2177 2273 2 2131 275 2057 OAI222S $T=594580 598200 1 180 $X=589000 $Y=597820
X3753 2110 2247 1 2253 2273 2 2295 282 2322 OAI222S $T=595820 618360 0 0 $X=595820 $Y=617980
X3754 2338 2141 1 2197 2273 2 2188 281 2057 OAI222S $T=603880 598200 1 180 $X=598300 $Y=597820
X3755 2110 2340 1 2296 2273 2 2328 287 2322 OAI222S $T=607600 618360 1 180 $X=602020 $Y=617980
X3756 2338 2173 1 2229 2273 2 2249 290 2345 OAI222S $T=613180 588120 1 180 $X=607600 $Y=587740
X3757 2369 2299 1 2267 2379 2 2334 2394 2391 OAI222S $T=612560 648600 1 0 $X=612560 $Y=643180
X3758 2369 2357 1 2309 2379 2 2378 2392 2391 OAI222S $T=613180 648600 0 0 $X=613180 $Y=648220
X3759 2338 2350 1 2390 2273 2 2349 297 2345 OAI222S $T=622480 598200 0 180 $X=616900 $Y=592780
X3760 2338 2331 1 2236 2406 2 2260 298 2322 OAI222S $T=624960 567960 1 180 $X=619380 $Y=567580
X3761 2410 2409 1 2354 1931 2 2415 2421 2402 OAI222S $T=626820 688920 0 180 $X=621240 $Y=683500
X3762 2410 2384 1 2288 2379 2 2399 2418 2402 OAI222S $T=628060 658680 1 180 $X=622480 $Y=658300
X3763 2400 2303 1 2277 2406 2 2218 304 2431 OAI222S $T=626200 557880 1 0 $X=626200 $Y=552460
X3764 2369 2403 1 2438 2435 2 2412 2437 2391 OAI222S $T=632400 628440 0 180 $X=626820 $Y=623020
X3765 2338 2430 1 2372 2434 2 2411 306 2322 OAI222S $T=628060 578040 0 0 $X=628060 $Y=577660
X3766 2400 309 1 2248 2406 2 2191 305 2431 OAI222S $T=636120 547800 1 180 $X=630540 $Y=547420
X3767 2410 2464 1 2373 2448 2 2443 2451 2402 OAI222S $T=636120 658680 0 180 $X=630540 $Y=653260
X3768 2369 2476 1 2474 2435 2 2427 2468 2391 OAI222S $T=639840 628440 1 180 $X=634260 $Y=628060
X3769 2494 2487 1 2268 2448 2 2477 2483 2459 OAI222S $T=644800 658680 1 180 $X=639220 $Y=658300
X3770 2400 2478 1 2396 2434 2 2356 323 2431 OAI222S $T=642940 567960 1 0 $X=642940 $Y=562540
X3771 2369 2498 1 2503 2435 2 2502 2510 2391 OAI222S $T=648520 628440 1 180 $X=642940 $Y=628060
X3772 2400 2408 1 2355 2434 2 2432 324 2431 OAI222S $T=643560 557880 1 0 $X=643560 $Y=552460
X3773 2400 2501 1 2485 2434 2 2473 325 2431 OAI222S $T=643560 557880 0 0 $X=643560 $Y=557500
X3774 2494 2530 1 2300 2448 2 2511 2525 2459 OAI222S $T=653480 658680 1 180 $X=647900 $Y=658300
X3775 2494 2551 1 2194 2448 2 2522 2549 2459 OAI222S $T=657200 658680 0 180 $X=651620 $Y=653260
X3776 2494 2570 1 2256 2448 2 2543 2565 2459 OAI222S $T=660920 658680 1 180 $X=655340 $Y=658300
X3777 2494 2568 1 2535 2435 2 2550 2579 2459 OAI222S $T=665880 638520 0 180 $X=660300 $Y=633100
X3778 2494 2577 1 2556 2435 2 2540 2582 2459 OAI222S $T=666500 628440 1 180 $X=660920 $Y=628060
X3779 1794 116 1679 2 1 167 170 116 165 180 675 ICV_12 $T=482980 547800 1 0 $X=482980 $Y=542380
X3780 1800 116 165 2 1 1884 1888 116 165 1930 675 ICV_12 $T=484220 547800 0 0 $X=484220 $Y=547420
X3781 2024 1791 2009 2 1 2074 2079 1791 2052 2117 675 ICV_12 $T=528240 668760 1 0 $X=528240 $Y=663340
X3782 2061 152 2108 2 1 2077 2120 152 2108 2158 675 ICV_12 $T=540640 699000 1 0 $X=540640 $Y=693580
X3783 2171 1791 2148 2 1 2201 1845 1791 2237 2262 675 ICV_12 $T=564820 608280 0 0 $X=564820 $Y=607900
X3784 2180 250 260 2 1 2209 2224 250 273 2255 675 ICV_12 $T=566680 547800 0 0 $X=566680 $Y=547420
X3785 2181 1791 2207 2 1 2220 2228 1791 2207 2271 675 ICV_12 $T=567300 648600 0 0 $X=567300 $Y=648220
X3786 1849 1791 2237 2 1 2278 2284 2290 2237 2332 675 ICV_12 $T=580320 598200 1 0 $X=580320 $Y=592780
X3787 2234 1791 2266 2 1 2276 2291 2290 2266 2315 675 ICV_12 $T=581560 628440 0 0 $X=581560 $Y=628060
X3788 312 271 2505 2 1 2508 326 271 2505 2538 675 ICV_12 $T=636120 719160 1 0 $X=636120 $Y=713740
X3789 2555 271 2462 2 1 2581 337 271 2611 349 675 ICV_12 $T=655340 678840 1 0 $X=655340 $Y=673420
X3790 2572 2290 2600 2 1 2596 2394 2290 2621 2649 675 ICV_12 $T=663400 638520 0 0 $X=663400 $Y=638140
X3791 2579 2290 2621 2 1 2630 2510 2290 2668 2685 675 ICV_12 $T=670840 638520 1 0 $X=670840 $Y=633100
X3792 2483 2290 2618 2 1 2656 2525 2290 2668 2719 675 ICV_12 $T=677040 648600 0 0 $X=677040 $Y=648220
X3793 1818 439 457 2 1 3531 464 439 469 3578 675 ICV_12 $T=810960 547800 1 0 $X=810960 $Y=542380
X3794 482 465 3547 2 1 3628 3518 465 3637 3713 675 ICV_12 $T=838860 648600 0 0 $X=838860 $Y=648220
X3795 4281 4080 4309 2 1 4320 4320 4080 4313 4354 675 ICV_12 $T=968440 628440 0 0 $X=968440 $Y=628060
X3796 4365 624 4387 2 1 4398 4398 624 4387 4424 675 ICV_12 $T=994480 678840 0 0 $X=994480 $Y=678460
X3797 4408 4080 4410 2 1 4412 4436 4080 4455 4460 675 ICV_12 $T=1009360 618360 0 0 $X=1009360 $Y=617980
X3798 646 585 644 2 1 4480 4480 585 644 651 675 ICV_12 $T=1028580 547800 1 0 $X=1028580 $Y=542380
X3799 867 2 1 851 BUF3 $T=316820 638520 1 0 $X=316820 $Y=633100
X3800 1121 2 1 1147 BUF3 $T=355880 638520 0 0 $X=355880 $Y=638140
X3801 976 2 1 1382 BUF3 $T=393080 638520 0 0 $X=393080 $Y=638140
X3802 1389 2 1 1165 BUF3 $T=396800 648600 0 180 $X=393080 $Y=643180
X3803 111 2 1 122 BUF3 $T=437100 709080 0 0 $X=437100 $Y=708700
X3804 175 2 1 1764 BUF3 $T=506540 699000 0 180 $X=502820 $Y=693580
X3805 2052 2 1 2067 BUF3 $T=537540 648600 1 0 $X=537540 $Y=643180
X3806 2067 2 1 2002 BUF3 $T=538780 628440 0 0 $X=538780 $Y=628060
X3807 2123 2 1 260 BUF3 $T=572880 578040 1 0 $X=572880 $Y=572620
X3808 633 2 1 631 BUF3 $T=1001920 688920 0 180 $X=998200 $Y=683500
X3809 4551 2 1 4510 BUF3 $T=1070120 598200 1 180 $X=1066400 $Y=597820
X3810 4601 2 1 658 BUF3 $T=1116620 557880 1 180 $X=1112900 $Y=557500
X3811 2002 1971 1 2 INV6 $T=522040 618360 1 180 $X=517080 $Y=617980
X3812 1566 1 1453 2 BUF4CK $T=434620 648600 0 180 $X=429660 $Y=643180
X3813 1858 1 1865 2 BUF4CK $T=501580 638520 0 0 $X=501580 $Y=638140
X3814 1895 1 1894 2 BUF4CK $T=506540 648600 1 0 $X=506540 $Y=643180
X3815 2096 1 1963 2 BUF4CK $T=546840 578040 1 180 $X=541880 $Y=577660
X3816 2110 1 1927 2 BUF4CK $T=548700 588120 0 180 $X=543740 $Y=582700
X3817 2627 1 2628 2 BUF4CK $T=683860 618360 1 0 $X=683860 $Y=612940
X3818 2703 1 2718 2 BUF4CK $T=701220 608280 1 0 $X=701220 $Y=602860
X3819 2758 1 2682 2 BUF4CK $T=709900 628440 0 0 $X=709900 $Y=628060
X3820 2069 184 1 2 INV8CK $T=538780 688920 0 0 $X=538780 $Y=688540
X3821 523 524 1 2 INV8CK $T=881020 557880 0 0 $X=881020 $Y=557500
X3822 679 690 1 2 INV4CK $T=262260 618360 1 0 $X=262260 $Y=612940
X3823 1955 216 1 2 INV4CK $T=531340 547800 0 0 $X=531340 $Y=547420
X3824 2286 2069 1 2 INV4CK $T=592720 688920 0 0 $X=592720 $Y=688540
X3825 523 4324 1 2 INV4CK $T=980220 547800 0 0 $X=980220 $Y=547420
X3826 906 904 896 2 1 928 XOR3 $T=314960 678840 1 0 $X=314960 $Y=673420
X3827 3092 3245 3269 2 1 3304 XOR3 $T=776860 578040 0 0 $X=776860 $Y=577660
X3828 3253 3165 3256 2 1 3408 XOR3 $T=790500 678840 0 0 $X=790500 $Y=678460
X3829 728 722 734 683 1 2 ND3P $T=275900 608280 0 180 $X=270940 $Y=602860
X3830 728 720 742 708 1 2 ND3P $T=277140 578040 1 180 $X=272180 $Y=577660
X3831 722 712 691 717 1 2 ND3P $T=272800 608280 0 0 $X=272800 $Y=607900
X3832 728 748 742 752 1 2 ND3P $T=283960 588120 0 180 $X=279000 $Y=582700
X3833 742 822 728 776 1 2 ND3P $T=288920 578040 0 0 $X=288920 $Y=577660
X3834 811 800 794 742 1 2 ND3P $T=296980 588120 0 180 $X=292020 $Y=582700
X3835 822 843 819 804 1 2 ND3P $T=294500 578040 1 0 $X=294500 $Y=572620
X3836 880 811 885 862 1 2 ND3P $T=310000 588120 1 0 $X=310000 $Y=582700
X3837 1602 1585 1599 1613 1 2 ND3P $T=438340 678840 1 0 $X=438340 $Y=673420
X3838 3293 3247 3309 3282 1 2 ND3P $T=786160 658680 1 180 $X=781200 $Y=658300
X3839 3356 3293 3331 3370 1 2 ND3P $T=791740 658680 0 0 $X=791740 $Y=658300
X3840 3426 3406 3446 3412 1 2 ND3P $T=806620 598200 1 180 $X=801660 $Y=597820
X3841 3483 3498 3491 3492 1 2 ND3P $T=810960 598200 0 0 $X=810960 $Y=597820
X3842 456 3503 3505 3504 1 2 ND3P $T=815300 699000 1 0 $X=815300 $Y=693580
X3843 3524 3509 3535 3511 1 2 ND3P $T=824600 608280 1 180 $X=819640 $Y=607900
X3844 3351 3523 3527 3401 1 2 ND3P $T=825220 668760 1 180 $X=820260 $Y=668380
X3845 3523 3572 3515 3345 1 2 ND3P $T=827700 668760 0 0 $X=827700 $Y=668380
X3846 3742 3775 3785 3771 1 2 ND3P $T=877920 699000 1 180 $X=872960 $Y=698620
X3847 4249 4286 4129 4287 1 2 ND3P $T=974020 688920 1 180 $X=969060 $Y=688540
X3848 4129 4293 4249 4300 1 2 ND3P $T=976500 688920 0 180 $X=971540 $Y=683500
X3849 4286 4290 4307 4308 1 2 ND3P $T=972780 699000 0 0 $X=972780 $Y=698620
X3850 700 731 683 1 2 OR2P $T=275900 658680 0 180 $X=272180 $Y=653260
X3851 2876 2860 380 1 2 OR2P $T=727260 547800 0 180 $X=723540 $Y=542380
X3852 3279 3180 3301 1 2 OR2P $T=781200 648600 0 0 $X=781200 $Y=648220
X3853 3236 3327 3401 1 2 OR2P $T=795460 668760 0 0 $X=795460 $Y=668380
X3854 3339 3365 3424 1 2 OR2P $T=797320 567960 1 0 $X=797320 $Y=562540
X3855 3418 3449 3510 1 2 OR2P $T=820260 638520 1 0 $X=820260 $Y=633100
X3856 4196 4190 4207 1 2 OR2P $T=944260 699000 1 0 $X=944260 $Y=693580
X3857 750 2 1 676 742 NR2F $T=279620 598200 1 180 $X=272800 $Y=597820
X3858 783 2 1 809 684 NR2F $T=288300 608280 1 0 $X=288300 $Y=602860
X3859 1225 2 1 1199 1154 NR2F $T=366420 699000 1 180 $X=359600 $Y=698620
X3860 3482 2 1 3474 3370 NR2F $T=811580 668760 1 0 $X=811580 $Y=663340
X3861 4207 2 1 4238 4249 NR2F $T=961000 688920 1 180 $X=954180 $Y=688540
X3862 711 3 738 749 4639 1 2 DFFRBP $T=267220 557880 1 0 $X=267220 $Y=552460
X3863 744 3 738 4 4640 1 2 DFFRBP $T=277140 547800 0 0 $X=277140 $Y=547420
X3864 39 11 942 4641 982 1 2 DFFRBP $T=339760 699000 0 180 $X=325500 $Y=693580
X3865 3262 465 3700 4642 3716 1 2 DFFRBP $T=849400 658680 1 0 $X=849400 $Y=653260
X3866 4215 4080 4185 4133 4036 1 2 DFFRBP $T=951080 668760 0 180 $X=936820 $Y=663340
X3867 4361 624 4333 4230 4643 1 2 DFFRBP $T=994480 668760 1 180 $X=980220 $Y=668380
X3868 2643 1 2 2659 INV3CK $T=688200 598200 1 0 $X=688200 $Y=592780
X3869 976 1018 1 2 INV12 $T=381300 648600 0 0 $X=381300 $Y=648220
X3870 1158 1128 1 1133 922 2 OAI12HP $T=358980 588120 0 180 $X=348440 $Y=582700
X3871 1181 1154 1 1144 1060 2 OAI12HP $T=363320 699000 0 180 $X=352780 $Y=693580
X3872 86 1494 1 1535 1335 2 OAI12HP $T=419120 709080 0 0 $X=419120 $Y=708700
X3873 3493 3479 1 3455 3391 2 OAI12HP $T=816540 628440 0 180 $X=806000 $Y=623020
X3874 4238 4218 1 4245 4264 2 OAI12HP $T=955420 699000 1 0 $X=955420 $Y=693580
X3875 15 11 7 815 1 2 4644 DFFRBN $T=306900 719160 0 180 $X=293880 $Y=713740
X3876 20 11 7 853 1 2 4645 DFFRBN $T=313100 709080 1 180 $X=300080 $Y=708700
X3877 1084 3 29 1052 1 2 1038 DFFRBN $T=349060 557880 0 180 $X=336040 $Y=552460
X3878 3590 465 3637 3662 1 2 4646 DFFRBN $T=837000 658680 0 0 $X=837000 $Y=658300
X3879 3540 465 3637 3703 1 2 4647 DFFRBN $T=847540 648600 1 0 $X=847540 $Y=643180
X3880 4089 4080 4047 3919 1 2 4648 DFFRBN $T=927520 668760 1 180 $X=914500 $Y=668380
X3881 4189 4080 4047 4056 1 2 4649 DFFRBN $T=941160 678840 0 180 $X=928140 $Y=673420
X3882 4267 4080 4239 4221 1 2 4650 DFFRBN $T=965340 668760 0 180 $X=952320 $Y=663340
X3883 807 1 832 800 2 841 ND3HT $T=301940 588120 1 180 $X=294500 $Y=587740
X3884 862 1 880 885 2 728 ND3HT $T=301940 588120 1 0 $X=301940 $Y=582700
X3885 916 1 959 971 2 880 ND3HT $T=317440 578040 0 0 $X=317440 $Y=577660
X3886 1034 1 30 986 2 26 ND3HT $T=333560 719160 0 180 $X=326120 $Y=713740
X3887 1034 1 30 986 2 37 ND3HT $T=333560 719160 1 0 $X=333560 $Y=713740
X3888 1039 1 1062 1071 2 986 ND3HT $T=336040 699000 0 0 $X=336040 $Y=698620
X3889 1279 1 1302 1305 2 971 ND3HT $T=375100 578040 0 0 $X=375100 $Y=577660
X3890 1324 1 1354 1361 2 1305 ND3HT $T=386260 578040 0 0 $X=386260 $Y=577660
X3891 1366 1 1379 1390 2 1071 ND3HT $T=391840 678840 0 0 $X=391840 $Y=678460
X3892 1467 1 1426 1487 2 1390 ND3HT $T=411680 678840 0 0 $X=411680 $Y=678460
X3893 1521 1 1508 1543 2 1502 ND3HT $T=422840 598200 0 0 $X=422840 $Y=597820
X3894 383 1 2817 380 2 386 ND3HT $T=722920 547800 0 180 $X=715480 $Y=542380
X3895 3370 1 3337 3351 2 3375 ND3HT $T=799180 658680 0 180 $X=791740 $Y=653260
X3896 3348 1 3326 3375 2 3354 ND3HT $T=792360 648600 1 0 $X=792360 $Y=643180
X3897 440 1 3315 444 2 3385 ND3HT $T=795460 547800 0 0 $X=795460 $Y=547420
X3898 3252 1 3416 3411 2 3427 ND3HT $T=807240 648600 0 180 $X=799800 $Y=643180
X3899 3370 1 3395 3351 2 3411 ND3HT $T=799800 658680 1 0 $X=799800 $Y=653260
X3900 440 1 3315 444 2 3454 ND3HT $T=810960 547800 0 180 $X=803520 $Y=542380
X3901 3496 1 3512 3503 2 3356 ND3HT $T=822740 688920 0 180 $X=815300 $Y=683500
X3902 3530 1 3480 3385 2 3524 ND3HT $T=823980 598200 0 180 $X=816540 $Y=592780
X3903 3798 1 3824 3775 2 3830 ND3HT $T=885980 699000 0 180 $X=878540 $Y=693580
X3904 4023 1 3970 3830 2 4016 ND3HT $T=915740 688920 0 180 $X=908300 $Y=683500
X3905 4079 1 4102 4016 2 4129 ND3HT $T=931860 688920 0 180 $X=924420 $Y=683500
X3906 4079 1 4102 4016 2 4162 ND3HT $T=939300 688920 0 180 $X=931860 $Y=683500
X3907 1191 1186 1150 1183 1 1177 2 AOI22S $T=363940 658680 1 180 $X=360220 $Y=658300
X3908 1187 1191 1049 1186 1 1177 2 AOI22S $T=366420 668760 1 180 $X=362700 $Y=668380
X3909 1249 1244 774 1241 1 1177 2 AOI22S $T=372620 668760 1 180 $X=368900 $Y=668380
X3910 1244 1186 958 1216 1 1177 2 AOI22S $T=371380 678840 1 0 $X=371380 $Y=673420
X3911 1183 1269 1195 1241 1 1177 2 AOI22S $T=373240 658680 0 0 $X=373240 $Y=658300
X3912 1369 1337 1332 1291 1 1241 2 AOI22S $T=390600 658680 0 180 $X=386880 $Y=653260
X3913 1428 1433 1439 1504 1 1471 2 AOI22S $T=418500 648600 0 0 $X=418500 $Y=648220
X3914 1538 1565 1561 1433 1 1471 2 AOI22S $T=432140 638520 1 0 $X=432140 $Y=633100
X3915 1608 1433 1601 1499 1 1471 2 AOI22S $T=441440 638520 1 180 $X=437720 $Y=638140
X3916 2653 2680 2706 2644 1 2657 2 AOI22S $T=696260 567960 1 180 $X=692540 $Y=567580
X3917 2698 2680 2700 2688 1 2657 2 AOI22S $T=696880 578040 1 0 $X=696880 $Y=572620
X3918 2787 2647 2782 2680 1 2736 2 AOI22S $T=711760 578040 0 180 $X=708040 $Y=572620
X3919 2974 2922 2942 2953 1 2736 2 AOI22S $T=734080 567960 1 180 $X=730360 $Y=567580
X3920 3019 2953 3009 2974 1 2736 2 AOI22S $T=740280 567960 1 180 $X=736560 $Y=567580
X3921 3041 2953 3063 3019 1 3045 2 AOI22S $T=748340 567960 1 180 $X=744620 $Y=567580
X3922 3078 2953 3123 3041 1 3045 2 AOI22S $T=759500 567960 1 180 $X=755780 $Y=567580
X3923 3126 2953 3133 3078 1 3045 2 AOI22S $T=759500 578040 0 180 $X=755780 $Y=572620
X3924 2962 2957 3114 3124 1 3045 2 AOI22S $T=755780 598200 1 0 $X=755780 $Y=592780
X3925 3062 425 3142 3121 1 2741 2 AOI22S $T=759500 688920 1 0 $X=759500 $Y=683500
X3926 3135 3126 3157 2957 1 3045 2 AOI22S $T=764460 588120 1 180 $X=760740 $Y=587740
X3927 3124 2957 3169 3135 1 3045 2 AOI22S $T=765080 598200 0 180 $X=761360 $Y=592780
X3928 3137 3118 3173 425 1 2741 2 AOI22S $T=766940 688920 1 180 $X=763220 $Y=688540
X3929 3118 3167 3183 425 1 427 2 AOI22S $T=766940 699000 0 180 $X=763220 $Y=693580
X3930 3167 428 3174 425 1 427 2 AOI22S $T=767560 709080 1 180 $X=763840 $Y=708700
X3931 3121 3137 3194 425 1 2741 2 AOI22S $T=768180 688920 0 180 $X=764460 $Y=683500
X3932 1499 1 2 1295 BUF1CK $T=419740 638520 0 180 $X=417260 $Y=633100
X3933 1880 1 2 1854 BUF1CK $T=497240 678840 0 0 $X=497240 $Y=678460
X3934 2057 1 2 2345 BUF1CK $T=609460 598200 1 0 $X=609460 $Y=592780
X3935 2618 1 2 2600 BUF1CK $T=680140 658680 0 180 $X=677660 $Y=653260
X3936 2611 1 2 2557 BUF1CK $T=683860 668760 1 180 $X=681380 $Y=668380
X3937 2369 1 2 2110 BUF8CK $T=616280 618360 1 180 $X=607600 $Y=617980
X3938 2402 1 2 2391 BUF8CK $T=627440 648600 1 180 $X=618760 $Y=648220
X3939 691 686 1 681 679 2 OAI12H $T=264740 618360 1 180 $X=258540 $Y=617980
X3940 755 753 1 743 716 2 OAI12H $T=282100 628440 0 180 $X=275900 $Y=623020
X3941 1050 1016 1 1030 789 2 OAI12H $T=337900 678840 1 180 $X=331700 $Y=678460
X3942 51 1157 1 1149 1107 2 OAI12H $T=358980 719160 0 180 $X=352780 $Y=713740
X3943 1217 52 1 54 1149 2 OAI12H $T=367660 719160 0 180 $X=361460 $Y=713740
X3944 1221 1165 1 1161 1190 2 OAI12H $T=368280 648600 0 180 $X=362080 $Y=643180
X3945 1312 1165 1 1296 1266 2 OAI12H $T=383160 648600 0 180 $X=376960 $Y=643180
X3946 1371 1017 1 976 1311 2 OAI12H $T=397420 618360 0 180 $X=391220 $Y=612940
X3947 1389 1473 1 1489 1484 2 OAI12H $T=422220 628440 1 180 $X=416020 $Y=628060
X3948 1572 1604 1 1582 1581 2 OAI12H $T=443300 608280 1 180 $X=437100 $Y=607900
X3949 1659 1653 1 1647 1636 2 OAI12H $T=453840 688920 0 180 $X=447640 $Y=683500
X3950 2634 2648 1 2654 2643 2 OAI12H $T=691920 598200 1 180 $X=685720 $Y=597820
X3951 2648 2634 1 2654 2701 2 OAI12H $T=691920 598200 0 0 $X=691920 $Y=597820
X3952 2682 2635 1 2690 2722 2 OAI12H $T=695020 618360 0 0 $X=695020 $Y=617980
X3953 2716 2664 1 2752 375 2 OAI12H $T=704320 547800 1 0 $X=704320 $Y=542380
X3954 2868 2877 1 2905 2916 2 OAI12H $T=721060 567960 1 0 $X=721060 $Y=562540
X3955 2941 2950 1 2908 2980 2 OAI12H $T=730360 547800 1 0 $X=730360 $Y=542380
X3956 3355 3346 1 3332 3399 2 OAI12H $T=792980 588120 1 0 $X=792980 $Y=582700
X3957 3466 3464 1 3488 3499 2 OAI12H $T=809100 699000 0 0 $X=809100 $Y=698620
X3958 3510 3492 1 3494 3478 2 OAI12H $T=819640 628440 1 180 $X=813440 $Y=628060
X3959 3714 501 1 3704 508 2 OAI12H $T=861800 567960 1 0 $X=861800 $Y=562540
X3960 3841 3836 1 3815 3867 2 OAI12H $T=884120 567960 0 0 $X=884120 $Y=567580
X3961 3892 3945 1 3944 3983 2 OAI12H $T=900860 688920 0 0 $X=900860 $Y=688540
X3962 618 4312 1 626 4369 2 OAI12H $T=988280 699000 0 0 $X=988280 $Y=698620
X3963 742 728 2 730 719 1 AOI12H $T=278380 588120 0 180 $X=272180 $Y=582700
X3964 734 728 2 758 760 1 AOI12H $T=279620 608280 1 0 $X=279620 $Y=602860
X3965 362 361 2 2664 359 1 AOI12H $T=693780 547800 0 180 $X=687580 $Y=542380
X3966 3456 3321 2 3484 3463 1 AOI12H $T=815920 648600 0 180 $X=809720 $Y=643180
X3967 3370 3351 2 3507 3321 1 AOI12H $T=810960 658680 1 0 $X=810960 $Y=653260
X3968 3480 3385 2 3513 3461 1 AOI12H $T=813440 588120 1 0 $X=813440 $Y=582700
X3969 3489 3351 2 3502 3465 1 AOI12H $T=819640 678840 0 180 $X=813440 $Y=673420
X3970 3527 3351 2 3548 3520 1 AOI12H $T=820880 658680 0 0 $X=820880 $Y=658300
X3971 1725 137 1734 1 2 1744 HA1 $T=461900 608280 1 0 $X=461900 $Y=602860
X3972 470 2262 3566 1 2 3555 HA1 $T=825840 608280 0 0 $X=825840 $Y=607900
X3973 3740 3765 3791 1 2 3806 HA1 $T=871100 588120 1 0 $X=871100 $Y=582700
X3974 3710 3739 3804 1 2 3835 HA1 $T=871720 567960 1 0 $X=871720 $Y=562540
X3975 3720 3779 3793 1 2 3821 HA1 $T=876680 578040 1 0 $X=876680 $Y=572620
X3976 3753 3855 3823 1 2 3816 HA1 $T=888460 588120 1 180 $X=880400 $Y=587740
X3977 3923 4017 4061 1 2 4078 HA1 $T=914500 567960 0 0 $X=914500 $Y=567580
X3978 3992 4025 4087 1 2 4075 HA1 $T=916980 557880 1 0 $X=916980 $Y=552460
X3979 3831 3979 4099 1 2 4082 HA1 $T=918840 598200 0 0 $X=918840 $Y=597820
X3980 1524 3 103 2 1 1577 1577 1588 675 ICV_17 $T=424080 547800 0 0 $X=424080 $Y=547420
X3981 1755 11 151 2 1 1817 1817 153 675 ICV_17 $T=470580 719160 1 0 $X=470580 $Y=713740
X3982 1833 1791 1842 2 1 1882 1881 1847 675 ICV_17 $T=483600 608280 1 0 $X=483600 $Y=602860
X3983 1862 1791 1896 2 1 1911 1911 1903 675 ICV_17 $T=491040 598200 1 0 $X=491040 $Y=592780
X3984 183 116 196 2 1 1994 1994 187 675 ICV_17 $T=509020 547800 1 0 $X=509020 $Y=542380
X3985 1953 116 1896 2 1 2008 2008 1906 675 ICV_17 $T=512120 598200 1 0 $X=512120 $Y=592780
X3986 2011 152 1986 2 1 2053 2053 219 675 ICV_17 $T=523900 699000 1 0 $X=523900 $Y=693580
X3987 2020 116 2046 2 1 2064 2064 1966 675 ICV_17 $T=526380 578040 1 0 $X=526380 $Y=572620
X3988 2121 152 2146 2 1 2167 2163 2176 675 ICV_17 $T=553660 668760 0 0 $X=553660 $Y=668380
X3989 2129 1791 2164 2 1 2179 2179 1958 675 ICV_17 $T=555520 598200 1 0 $X=555520 $Y=592780
X3990 2160 250 260 2 1 2203 2203 262 675 ICV_17 $T=561720 547800 1 0 $X=561720 $Y=542380
X3991 2166 250 260 2 1 2211 2211 203 675 ICV_17 $T=563580 567960 0 0 $X=563580 $Y=567580
X3992 2205 152 2226 2 1 2242 2242 2238 675 ICV_17 $T=572880 709080 1 0 $X=572880 $Y=703660
X3993 2305 2290 2293 2 1 2361 2361 2296 675 ICV_17 $T=600160 648600 0 0 $X=600160 $Y=648220
X3994 2370 2290 2360 2 1 2424 2424 2229 675 ICV_17 $T=613180 588120 1 0 $X=613180 $Y=582700
X3995 2407 2290 2360 2 1 2455 2455 2372 675 ICV_17 $T=620620 598200 0 0 $X=620620 $Y=597820
X3996 2519 2290 2589 2 1 2604 2588 2589 675 ICV_17 $T=661540 608280 1 0 $X=661540 $Y=602860
X3997 2560 2290 2600 2 1 2606 2606 2556 675 ICV_17 $T=662780 648600 1 0 $X=662780 $Y=643180
X3998 2564 2290 2600 2 1 2608 2608 2550 675 ICV_17 $T=663400 648600 0 0 $X=663400 $Y=648220
X3999 4460 4451 4474 2 1 4486 4471 4491 675 ICV_17 $T=1032920 618360 0 0 $X=1032920 $Y=617980
X4000 708 1 685 707 2 ND2T $T=265980 588120 0 180 $X=261020 $Y=582700
X4001 916 1 922 862 2 ND2T $T=310620 578040 0 0 $X=310620 $Y=577660
X4002 1060 1 1039 1034 2 ND2T $T=338520 709080 1 180 $X=333560 $Y=708700
X4003 1326 1 1311 1299 2 ND2T $T=385020 618360 0 180 $X=380060 $Y=612940
X4004 1480 1 1502 1361 2 ND2T $T=416020 598200 1 0 $X=416020 $Y=592780
X4005 86 1 1509 1535 2 ND2T $T=432140 709080 0 0 $X=432140 $Y=708700
X4006 3401 1 3433 3474 2 ND2T $T=810340 668760 0 180 $X=805380 $Y=663340
X4007 616 1 609 4318 2 ND2T $T=981460 709080 0 180 $X=976500 $Y=703660
X4008 60 63 1297 2 1 1331 XNR3 $T=374480 709080 1 0 $X=374480 $Y=703660
X4009 3154 3161 3223 2 1 3211 XNR3 $T=763220 567960 1 0 $X=763220 $Y=562540
X4010 3260 3212 3299 2 1 3323 XNR3 $T=778720 608280 1 0 $X=778720 $Y=602860
X4011 2856 3391 445 2879 1 2 MXL2H $T=796700 628440 1 0 $X=796700 $Y=623020
X4012 3396 3406 447 3453 1 2 MXL2H $T=799180 608280 1 0 $X=799180 $Y=602860
X4013 4280 4290 4215 4269 1 2 MXL2H $T=972780 699000 1 180 $X=964100 $Y=698620
X4014 1838 1 1883 2 BUF6CK $T=489800 668760 0 0 $X=489800 $Y=668380
X4015 1989 1 211 2 BUF6CK $T=522040 547800 1 0 $X=522040 $Y=542380
X4016 2057 1 1988 2 BUF6CK $T=535060 588120 0 0 $X=535060 $Y=587740
X4017 2410 1 2369 2 BUF6CK $T=626820 658680 0 180 $X=619380 $Y=653260
X4018 184 1555 1 2 INV6CK $T=509640 658680 0 0 $X=509640 $Y=658300
X4019 2351 2614 1 2 INV6CK $T=677660 658680 0 180 $X=672080 $Y=653260
X4020 4324 4394 1 2 INV6CK $T=1005640 598200 0 180 $X=1000060 $Y=592780
X4021 4324 4399 1 2 INV6CK $T=1013080 547800 0 180 $X=1007500 $Y=542380
X4022 1177 1216 2 1186 994 1187 1 AOI22H $T=368900 678840 0 180 $X=361460 $Y=673420
X4023 1291 1269 2 1186 1230 1337 1 AOI22H $T=380060 658680 0 0 $X=380060 $Y=658300
X4024 1417 1382 1389 1448 1 2 MXL2HP $T=401140 638520 0 0 $X=401140 $Y=638140
X4025 1883 1 2 1878 BUF3CK $T=510880 638520 1 180 $X=506540 $Y=638140
X4026 2110 1 2 2338 BUF3CK $T=611940 598200 1 0 $X=611940 $Y=592780
X4027 706 677 682 1 2 XNR2H $T=268460 638520 1 180 $X=259780 $Y=638140
X4028 694 714 741 1 2 XNR2H $T=262880 628440 0 0 $X=262880 $Y=628060
X4029 727 694 702 1 2 XNR2H $T=274660 638520 0 180 $X=265980 $Y=633100
X4030 770 727 747 1 2 XNR2H $T=287060 628440 1 180 $X=278380 $Y=628060
X4031 831 771 787 1 2 XNR2H $T=298840 618360 0 180 $X=290160 $Y=612940
X4032 817 770 795 1 2 XNR2H $T=300080 638520 0 180 $X=291400 $Y=633100
X4033 1217 1174 52 1 2 XNR2H $T=368900 709080 1 180 $X=360220 $Y=708700
X4034 1290 1287 1239 1 2 XNR2H $T=384400 588120 0 180 $X=375720 $Y=582700
X4035 3366 3336 3319 1 2 XNR2H $T=798560 578040 0 180 $X=789880 $Y=572620
X4036 2971 3373 3316 1 2 XNR2H $T=789880 608280 1 0 $X=789880 $Y=602860
X4037 3373 3363 3323 1 2 XNR2H $T=801040 598200 1 180 $X=792360 $Y=597820
X4038 960 1007 987 885 1 2 OA12P $T=329840 588120 0 180 $X=325500 $Y=582700
X4039 3180 3217 3185 3252 1 2 OA12P $T=773760 648600 1 0 $X=773760 $Y=643180
X4040 3254 3252 3229 3282 1 2 OA12P $T=777480 658680 1 0 $X=777480 $Y=653260
X4041 3402 3404 3390 3429 1 2 OA12P $T=801040 578040 0 0 $X=801040 $Y=577660
X4042 4026 4030 4070 4079 1 2 OA12P $T=918840 688920 0 0 $X=918840 $Y=688540
X4043 4196 4171 4211 4218 1 2 OA12P $T=949220 688920 0 0 $X=949220 $Y=688540
X4044 4251 4234 4250 4245 1 2 OA12P $T=962240 709080 0 180 $X=957900 $Y=703660
X4045 676 684 1 690 719 2 OAI12HT $T=254820 598200 0 0 $X=254820 $Y=597820
X4046 3474 3451 1 3403 3321 2 OAI12HT $T=815920 658680 1 180 $X=801040 $Y=658300
X4047 3436 3439 1 3429 3461 2 OAI12HT $T=803520 578040 1 0 $X=803520 $Y=572620
X4048 699 3 738 754 1 2 4651 DFFRBS $T=269080 557880 0 0 $X=269080 $Y=557500
X4049 821 3 738 766 1 2 4652 DFFRBS $T=296980 557880 0 180 $X=283960 $Y=552460
X4050 19 11 7 803 1 2 4653 DFFRBS $T=313100 699000 1 180 $X=300080 $Y=698620
X4051 24 11 7 908 1 2 4654 DFFRBS $T=323020 719160 0 180 $X=310000 $Y=713740
X4052 23 11 942 1006 1 2 4655 DFFRBS $T=320540 709080 1 0 $X=320540 $Y=703660
X4053 3389 465 3547 3641 1 2 4656 DFFRBS $T=833900 648600 1 0 $X=833900 $Y=643180
X4054 3470 465 3637 3701 1 2 4657 DFFRBS $T=846920 638520 0 0 $X=846920 $Y=638140
X4055 4265 4080 4185 4178 1 2 4658 DFFRBS $T=964720 668760 1 180 $X=951700 $Y=668380
X4056 4268 4080 4239 4170 1 2 4659 DFFRBS $T=965340 658680 1 180 $X=952320 $Y=658300
X4057 2142 250 2164 2 1 2187 2170 250 2123 2145 675 ICV_20 $T=571020 578040 0 180 $X=559240 $Y=572620
X4058 4045 4080 4205 2 1 4212 597 585 4182 4168 675 ICV_20 $T=950460 578040 0 180 $X=938680 $Y=572620
X4059 4276 4080 4247 2 1 4232 4233 4080 4247 4276 675 ICV_20 $T=955420 628440 1 0 $X=955420 $Y=623020
X4060 4246 4080 4213 2 1 4278 4278 4080 4041 4233 675 ICV_20 $T=969680 608280 0 180 $X=957900 $Y=602860
X4061 4337 585 4255 2 1 4272 4262 585 4330 4337 675 ICV_20 $T=975880 557880 1 0 $X=975880 $Y=552460
X4062 4378 585 4343 2 1 4344 4341 585 4330 4378 675 ICV_20 $T=989520 567960 1 0 $X=989520 $Y=562540
X4063 4400 624 4406 2 1 4430 4424 624 4406 4400 675 ICV_20 $T=1018040 688920 0 180 $X=1006260 $Y=683500
X4064 4432 4080 4437 2 1 4458 4457 4080 4437 4431 675 ICV_20 $T=1031680 638520 0 180 $X=1019900 $Y=633100
X4065 4435 624 4407 2 1 647 4397 624 4407 4434 675 ICV_20 $T=1032300 709080 0 180 $X=1020520 $Y=703660
X4066 4433 4080 4478 2 1 4492 4496 4451 4474 4464 675 ICV_20 $T=1046560 648600 0 180 $X=1034780 $Y=643180
X4067 4466 4451 4478 2 1 4494 4492 4451 4478 4466 675 ICV_20 $T=1047180 658680 0 180 $X=1035400 $Y=653260
X4068 4520 4451 4474 2 1 4495 4486 4451 4474 4530 675 ICV_20 $T=1049660 628440 1 0 $X=1049660 $Y=623020
X4069 4501 624 4509 2 1 4538 4516 624 4509 4501 675 ICV_20 $T=1061440 699000 0 180 $X=1049660 $Y=693580
X4070 4546 650 4532 2 1 4524 4524 650 4532 4563 675 ICV_20 $T=1061440 578040 1 0 $X=1061440 $Y=572620
X4071 4521 624 4517 2 1 4549 4547 624 4517 4521 675 ICV_20 $T=1073220 688920 0 180 $X=1061440 $Y=683500
X4072 4550 4451 4534 2 1 4515 4526 4451 4534 4550 675 ICV_20 $T=1062680 618360 1 0 $X=1062680 $Y=612940
X4073 4567 624 4514 2 1 4539 4539 4451 4562 4561 675 ICV_20 $T=1067640 668760 1 0 $X=1067640 $Y=663340
X4074 4558 650 4568 2 1 4578 4575 650 4568 4558 675 ICV_20 $T=1086860 588120 0 180 $X=1075080 $Y=582700
X4075 4578 4451 4551 2 1 4559 4560 650 4551 4575 675 ICV_20 $T=1075080 598200 1 0 $X=1075080 $Y=592780
X4076 4603 624 4566 2 1 4581 4584 624 4566 4603 675 ICV_20 $T=1088720 688920 1 0 $X=1088720 $Y=683500
X4077 4607 624 4562 2 1 4584 4586 624 4562 4607 675 ICV_20 $T=1089340 678840 1 0 $X=1089340 $Y=673420
X4078 4590 4451 4594 2 1 4609 4609 4451 4594 4583 675 ICV_20 $T=1101740 648600 0 180 $X=1089960 $Y=643180
X4079 4626 4451 4594 2 1 4611 4612 4451 4594 4626 675 ICV_20 $T=1103600 658680 1 0 $X=1103600 $Y=653260
X4080 4325 587 2 4063 1 620 MUX2S $T=981460 608280 1 0 $X=981460 $Y=602860
X4081 4349 587 2 4045 1 627 MUX2S $T=989520 598200 0 0 $X=989520 $Y=597820
X4082 4356 587 2 4058 1 630 MUX2S $T=992000 598200 1 0 $X=992000 $Y=592780
X4083 4373 632 2 3960 1 636 MUX2S $T=999440 588120 0 0 $X=999440 $Y=587740
X4084 4188 587 2 1 579 581 MUX2 $T=939300 598200 1 180 $X=934960 $Y=597820
X4085 4164 596 2 1 4194 4167 MUX2 $T=948600 557880 0 180 $X=944260 $Y=552460
X4086 4220 605 2 1 4223 4224 MUX2 $T=958520 557880 1 180 $X=954180 $Y=557500
X4087 4272 596 2 1 4294 4262 MUX2 $T=967820 557880 1 0 $X=967820 $Y=552460
X4088 615 613 2 1 4316 4283 MUX2 $T=974020 547800 0 0 $X=974020 $Y=547420
X4089 3441 3465 2 3451 3475 1 AOI12HP $T=802900 668760 0 0 $X=802900 $Y=668380
X4090 3450 3454 2 3479 3461 1 AOI12HP $T=804760 588120 0 0 $X=804760 $Y=587740
X4091 3653 3685 2 498 3645 1 AOI12HP $T=859940 567960 0 180 $X=849400 $Y=562540
X4092 616 4296 2 4312 4301 1 AOI12HP $T=982700 709080 1 180 $X=972160 $Y=708700
X4093 3621 3675 3647 3685 1 2 AO12P $T=850020 588120 0 0 $X=850020 $Y=587740
X4094 1297 63 1277 1217 1 2 MAO222P $T=377580 719160 1 0 $X=377580 $Y=713740
X4095 3270 3107 3224 3316 1 2 MAO222P $T=781200 598200 1 0 $X=781200 $Y=592780
X4096 2673 2671 2688 2 1 2681 AN3 $T=697500 588120 0 180 $X=693780 $Y=582700
X4097 1860 1865 1 1878 1877 1894 1723 1875 2 OAI222H $T=490420 638520 0 0 $X=490420 $Y=638140
X4098 1865 1972 1 1974 1878 1894 1739 2013 2 OAI222H $T=514600 638520 1 0 $X=514600 $Y=633100
X4099 234 237 1 2062 241 244 245 2073 2 OAI222H $T=541880 547800 1 0 $X=541880 $Y=542380
X4100 2073 2085 1 247 234 244 252 2124 2 OAI222H $T=566680 547800 1 180 $X=555520 $Y=547420
X4101 2400 267 1 288 2406 2431 302 285 2 OAI222H $T=619380 547800 0 0 $X=619380 $Y=547420
X4102 1389 1382 1513 1510 2 1 1526 MAOI1 $T=420360 638520 0 0 $X=420360 $Y=638140
X4103 1344 1018 1 2 BUF8 $T=388740 648600 0 0 $X=388740 $Y=648220
X4104 1174 1225 54 1 2 XNR2HP $T=357120 709080 1 0 $X=357120 $Y=703660
X4105 961 993 1 2 INV2CK $T=355260 608280 0 0 $X=355260 $Y=607900
X4106 683 680 2 676 1 ND2F $T=262260 608280 0 180 $X=256060 $Y=602860
.ENDS
***************************************
.SUBCKT ICV_22 1 2 3 4 5 6 7 8 9 10 11
** N=11 EP=11 IP=14 FDC=0
X0 1 2 3 4 5 6 QDFFRBN $T=0 0 0 0 $X=0 $Y=-380
X1 7 8 9 4 5 10 QDFFRBN $T=11780 10080 0 180 $X=0 $Y=4660
.ENDS
***************************************
.SUBCKT ICV_23 1 2 3 4 5 6 7 8 9 10 11
** N=11 EP=11 IP=14 FDC=0
X0 1 2 3 4 5 6 QDFFRBN $T=0 0 0 0 $X=0 $Y=-380
X1 7 8 9 4 5 10 QDFFRBN $T=12400 0 0 180 $X=620 $Y=-5420
.ENDS
***************************************
.SUBCKT OR2B1S I1 B1 GND O VCC
** N=6 EP=5 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT DFFRBT D CK RB Q GND VCC QB
** N=8 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT QDFFRBT D CK RB GND VCC Q
** N=7 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT INV1CK O I GND VCC
** N=5 EP=4 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT BUF2CK I O GND VCC
** N=5 EP=4 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MAOI1HP B1 B2 A2 A1 VCC GND O
** N=8 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OAI22HP B2 B1 GND A2 O A1 VCC
** N=8 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MOAI1HP B2 B1 GND A1 O A2 VCC
** N=8 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_24 1 2 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21
+ 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41
+ 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61
+ 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81
+ 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101
+ 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121
+ 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140 141
+ 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161
+ 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180 181
+ 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200 201
+ 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220 221
+ 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240 241
+ 242 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 259 260 261
+ 262 263 264 265 266 267 268 269 270 271 272 273 274 275 276 277 278 279 280 281
+ 282 283 284 285 286 287 288 289 290 291 292 293 294 295 296 297 298 299 300 301
+ 302 303 304 305 306 307 308 309 310 311 312 313 314 315 316 317 318 319 320 321
+ 322 323 324 325 326 327 328 329 330 331 332 333 334 335 336 337 338 339 340 341
+ 342 343 344 345 346 347 348 349 350 351 352 353 354 355 356 357 358 359 360 361
+ 362 363 364 365 366 367 368 369 370 371 372 373 374 375 376 377 378 379 380 381
+ 382 383 384 385 386 387 388 389 390 391 392 393 394 395 396 397 398 399 400 401
+ 402 403 404 405 406 407 408 409 410 411 412 413 414 415 416 417 418 419 420 421
+ 422 423 424 425 426 427 428 429 430 431 432 433 434 435 436 437 438 439 440 441
+ 442 443 444 445 446 447 448 449 450 451 452 453 454 455 456 457 458 459 460 461
+ 462 463 464 465 466 467 468 469 470 471 472 473 474 475 476 477 478 479 480 481
+ 482 483 484 485 486 487 488 489 490 491 492 493 494 495 496 497 498 499 500 501
+ 506
** N=3517 EP=501 IP=19511 FDC=0
X0 1165 1 2 1055 BUF1S $T=466240 416760 0 180 $X=463760 $Y=411340
X1 1516 1 2 1519 BUF1S $T=566680 436920 0 0 $X=566680 $Y=436540
X2 2621 1 2 2573 BUF1S $T=824600 477240 1 180 $X=822120 $Y=476860
X3 376 1 2 2766 BUF1S $T=868000 537720 1 0 $X=868000 $Y=532300
X4 2958 1 2 2863 BUF1S $T=911400 426840 0 180 $X=908920 $Y=421420
X5 2958 1 2 3210 BUF1S $T=987040 426840 0 180 $X=984560 $Y=421420
X6 462 1 2 2857 BUF1S $T=998820 447000 1 180 $X=996340 $Y=446620
X7 3253 1 2 463 BUF1S $T=1001920 537720 0 180 $X=999440 $Y=532300
X8 3210 1 2 3253 BUF1S $T=1000060 467160 0 0 $X=1000060 $Y=466780
X9 24 2 1 509 BUF1 $T=324880 527640 0 180 $X=322400 $Y=522220
X10 567 2 1 564 BUF1 $T=326740 477240 0 0 $X=326740 $Y=476860
X11 24 2 1 608 BUF1 $T=341000 527640 0 0 $X=341000 $Y=527260
X12 633 2 1 684 BUF1 $T=371380 436920 1 0 $X=371380 $Y=431500
X13 811 2 1 756 BUF1 $T=383780 467160 0 180 $X=381300 $Y=461740
X14 890 2 1 901 BUF1 $T=398040 517560 0 0 $X=398040 $Y=517180
X15 944 2 1 885 BUF1 $T=411060 477240 0 180 $X=408580 $Y=471820
X16 936 2 1 953 BUF1 $T=415400 457080 0 180 $X=412920 $Y=451660
X17 936 2 1 921 BUF1 $T=417260 487320 0 180 $X=414780 $Y=481900
X18 958 2 1 967 BUF1 $T=418500 507480 1 0 $X=418500 $Y=502060
X19 865 2 1 1057 BUF1 $T=436480 477240 0 0 $X=436480 $Y=476860
X20 925 2 1 1061 BUF1 $T=437720 457080 0 0 $X=437720 $Y=456700
X21 65 2 1 944 BUF1 $T=440200 497400 1 0 $X=440200 $Y=491980
X22 978 2 1 1082 BUF1 $T=440820 527640 0 0 $X=440820 $Y=527260
X23 1047 2 1 811 BUF1 $T=443300 457080 0 0 $X=443300 $Y=456700
X24 1132 2 1 979 BUF1 $T=453220 416760 1 180 $X=450740 $Y=416380
X25 1082 2 1 1125 BUF1 $T=450740 527640 1 0 $X=450740 $Y=522220
X26 949 2 1 1050 BUF1 $T=466240 426840 0 0 $X=466240 $Y=426460
X27 1194 2 1 82 BUF1 $T=469340 537720 0 180 $X=466860 $Y=532300
X28 1050 2 1 1202 BUF1 $T=467480 416760 0 0 $X=467480 $Y=416380
X29 1202 2 1 70 BUF1 $T=469960 406680 0 0 $X=469960 $Y=406300
X30 1233 2 1 1132 BUF1 $T=479880 416760 0 180 $X=477400 $Y=411340
X31 1253 2 1 1212 BUF1 $T=481740 507480 0 180 $X=479260 $Y=502060
X32 1202 2 1 1267 BUF1 $T=486700 416760 0 0 $X=486700 $Y=416380
X33 1280 2 1 1233 BUF1 $T=494760 426840 0 180 $X=492280 $Y=421420
X34 1267 2 1 1293 BUF1 $T=498480 447000 1 0 $X=498480 $Y=441580
X35 1309 2 1 1280 BUF1 $T=507160 457080 0 180 $X=504680 $Y=451660
X36 1267 2 1 1298 BUF1 $T=505920 426840 1 0 $X=505920 $Y=421420
X37 1305 2 1 1309 BUF1 $T=505920 477240 0 0 $X=505920 $Y=476860
X38 1305 2 1 1297 BUF1 $T=512120 517560 1 0 $X=512120 $Y=512140
X39 1297 2 1 113 BUF1 $T=513360 527640 0 0 $X=513360 $Y=527260
X40 1236 2 1 120 BUF1 $T=522040 517560 1 0 $X=522040 $Y=512140
X41 1375 2 1 1409 BUF1 $T=535060 457080 1 0 $X=535060 $Y=451660
X42 1417 2 1 1467 BUF1 $T=551180 517560 1 0 $X=551180 $Y=512140
X43 1483 2 1 1479 BUF1 $T=561720 447000 1 0 $X=561720 $Y=441580
X44 1524 2 1 1535 BUF1 $T=567920 447000 1 0 $X=567920 $Y=441580
X45 1543 2 1 1550 BUF1 $T=574740 436920 0 0 $X=574740 $Y=436540
X46 1563 2 1 1413 BUF1 $T=575360 527640 1 0 $X=575360 $Y=522220
X47 1556 2 1 1582 BUF1 $T=581560 477240 1 0 $X=581560 $Y=471820
X48 1525 2 1 173 BUF1 $T=582800 537720 1 0 $X=582800 $Y=532300
X49 1602 2 1 1619 BUF1 $T=588380 507480 1 0 $X=588380 $Y=502060
X50 1605 2 1 1574 BUF1 $T=594580 436920 1 180 $X=592100 $Y=436540
X51 187 2 1 1762 BUF1 $T=626820 537720 1 0 $X=626820 $Y=532300
X52 187 2 1 192 BUF1 $T=631780 537720 0 0 $X=631780 $Y=537340
X53 1835 2 1 1855 BUF1 $T=648520 477240 1 0 $X=648520 $Y=471820
X54 1889 2 1 223 BUF1 $T=662780 406680 1 0 $X=662780 $Y=401260
X55 1896 2 1 1888 BUF1 $T=675800 467160 1 180 $X=673320 $Y=466780
X56 234 2 1 242 BUF1 $T=675180 396600 1 0 $X=675180 $Y=391180
X57 1934 2 1 1925 BUF1 $T=682620 406680 0 180 $X=680140 $Y=401260
X58 1952 2 1 1953 BUF1 $T=683240 487320 0 0 $X=683240 $Y=486940
X59 240 2 1 1987 BUF1 $T=685100 527640 1 0 $X=685100 $Y=522220
X60 1892 2 1 1993 BUF1 $T=687580 507480 1 0 $X=687580 $Y=502060
X61 1940 2 1 259 BUF1 $T=689440 436920 0 0 $X=689440 $Y=436540
X62 2031 2 1 265 BUF1 $T=702460 406680 1 180 $X=699980 $Y=406300
X63 2057 2 1 2042 BUF1 $T=701840 477240 0 0 $X=701840 $Y=476860
X64 2038 2 1 269 BUF1 $T=702460 416760 1 0 $X=702460 $Y=411340
X65 1994 2 1 273 BUF1 $T=711760 426840 0 0 $X=711760 $Y=426460
X66 2125 2 1 2054 BUF1 $T=716100 467160 1 180 $X=713620 $Y=466780
X67 1993 2 1 2122 BUF1 $T=716100 517560 0 180 $X=713620 $Y=512140
X68 2107 2 1 2174 BUF1 $T=720440 436920 1 0 $X=720440 $Y=431500
X69 2520 2 1 2576 BUF1 $T=819640 507480 0 180 $X=817160 $Y=502060
X70 2560 2 1 337 BUF1 $T=820880 527640 1 180 $X=818400 $Y=527260
X71 2560 2 1 2679 BUF1 $T=827080 517560 0 0 $X=827080 $Y=517180
X72 2679 2 1 2670 BUF1 $T=832660 517560 0 0 $X=832660 $Y=517180
X73 2469 2 1 2717 BUF1 $T=844440 426840 0 0 $X=844440 $Y=426460
X74 2717 2 1 2731 BUF1 $T=849400 426840 0 0 $X=849400 $Y=426460
X75 2712 2 1 2706 BUF1 $T=856840 467160 0 0 $X=856840 $Y=466780
X76 2754 2 1 2712 BUF1 $T=860560 457080 1 180 $X=858080 $Y=456700
X77 2717 2 1 2754 BUF1 $T=858700 436920 0 0 $X=858700 $Y=436540
X78 2754 2 1 2784 BUF1 $T=863040 436920 0 0 $X=863040 $Y=436540
X79 2754 2 1 2785 BUF1 $T=863040 457080 0 0 $X=863040 $Y=456700
X80 2784 2 1 2770 BUF1 $T=872960 426840 1 180 $X=870480 $Y=426460
X81 2785 2 1 2877 BUF1 $T=888460 477240 1 0 $X=888460 $Y=471820
X82 2950 2 1 2909 BUF1 $T=910780 457080 1 0 $X=910780 $Y=451660
X83 2950 2 1 2986 BUF1 $T=922560 447000 0 0 $X=922560 $Y=446620
X84 3051 2 1 3052 BUF1 $T=931860 477240 0 0 $X=931860 $Y=476860
X85 429 2 1 417 BUF1 $T=937440 396600 0 180 $X=934960 $Y=391180
X86 2986 2 1 3051 BUF1 $T=934960 447000 0 0 $X=934960 $Y=446620
X87 3034 2 1 3063 BUF1 $T=936200 426840 0 0 $X=936200 $Y=426460
X88 3003 2 1 3075 BUF1 $T=938680 406680 0 0 $X=938680 $Y=406300
X89 3063 2 1 3079 BUF1 $T=941160 436920 1 0 $X=941160 $Y=431500
X90 3163 2 1 3134 BUF1 $T=964720 436920 0 180 $X=962240 $Y=431500
X91 3161 2 1 3164 BUF1 $T=977120 406680 1 180 $X=974640 $Y=406300
X92 451 2 1 3169 BUF1 $T=983320 527640 1 180 $X=980840 $Y=527260
X93 3171 2 1 3224 BUF1 $T=983320 477240 0 0 $X=983320 $Y=476860
X94 3173 2 1 3192 BUF1 $T=987660 447000 0 0 $X=987660 $Y=446620
X95 3224 2 1 3211 BUF1 $T=990140 477240 1 180 $X=987660 $Y=476860
X96 474 2 1 3250 BUF1 $T=1018040 507480 0 180 $X=1015560 $Y=502060
X97 3250 2 1 3292 BUF1 $T=1019900 507480 1 0 $X=1019900 $Y=502060
X98 3290 2 1 3294 BUF1 $T=1034160 477240 1 180 $X=1031680 $Y=476860
X99 474 2 1 3330 BUF1 $T=1039740 436920 0 0 $X=1039740 $Y=436540
X100 3330 2 1 3315 BUF1 $T=1050280 426840 1 180 $X=1047800 $Y=426460
X101 482 2 1 3396 BUF1 $T=1073220 537720 1 0 $X=1073220 $Y=532300
X102 489 2 1 490 BUF1 $T=1076320 416760 0 0 $X=1076320 $Y=416380
X103 3393 2 1 3401 BUF1 $T=1076320 447000 1 0 $X=1076320 $Y=441580
X104 3419 2 1 3417 BUF1 $T=1084380 416760 1 0 $X=1084380 $Y=411340
X105 3419 2 1 3440 BUF1 $T=1101120 416760 0 0 $X=1101120 $Y=416380
X106 500 2 1 501 BUF1 $T=1126540 467160 0 0 $X=1126540 $Y=466780
X107 510 8 509 2 1 507 QDFFRBN $T=300700 527640 0 180 $X=288920 $Y=522220
X108 533 8 509 2 1 15 QDFFRBN $T=319920 527640 1 180 $X=308140 $Y=527260
X109 590 8 24 2 1 22 QDFFRBN $T=336660 527640 1 180 $X=324880 $Y=527260
X110 649 8 608 2 1 30 QDFFRBN $T=352160 537720 0 180 $X=340380 $Y=532300
X111 664 8 608 2 1 34 QDFFRBN $T=358980 527640 1 180 $X=347200 $Y=527260
X112 48 8 45 2 1 49 QDFFRBN $T=398660 537720 0 0 $X=398660 $Y=537340
X113 50 8 55 2 1 58 QDFFRBN $T=412920 537720 0 0 $X=412920 $Y=537340
X114 1019 61 949 2 1 988 QDFFRBN $T=433380 416760 0 180 $X=421600 $Y=411340
X115 987 8 978 2 1 1015 QDFFRBN $T=424080 537720 1 0 $X=424080 $Y=532300
X116 1068 66 978 2 1 1034 QDFFRBN $T=445160 517560 1 180 $X=433380 $Y=517180
X117 1046 66 1082 2 1 1087 QDFFRBN $T=437100 537720 1 0 $X=437100 $Y=532300
X118 1083 61 70 2 1 1143 QDFFRBN $T=445160 396600 0 0 $X=445160 $Y=396220
X119 1089 61 70 2 1 1135 QDFFRBN $T=445780 406680 1 0 $X=445780 $Y=401260
X120 1091 66 1125 2 1 75 QDFFRBN $T=445780 527640 0 0 $X=445780 $Y=527260
X121 1097 66 1125 2 1 77 QDFFRBN $T=447020 517560 0 0 $X=447020 $Y=517180
X122 1144 61 1050 2 1 1092 QDFFRBN $T=459420 426840 0 180 $X=447640 $Y=421420
X123 1092 61 1050 2 1 1072 QDFFRBN $T=459420 426840 1 180 $X=447640 $Y=426460
X124 1099 66 1082 2 1 1159 QDFFRBN $T=449500 537720 1 0 $X=449500 $Y=532300
X125 1138 61 70 2 1 1196 QDFFRBN $T=455700 406680 0 0 $X=455700 $Y=406300
X126 1156 66 1082 2 1 73 QDFFRBN $T=467480 527640 0 180 $X=455700 $Y=522220
X127 1185 66 1082 2 1 76 QDFFRBN $T=469340 527640 1 180 $X=457560 $Y=527260
X128 1161 61 1050 2 1 1211 QDFFRBN $T=460660 426840 1 0 $X=460660 $Y=421420
X129 1238 66 1212 2 1 899 QDFFRBN $T=480500 527640 0 180 $X=468720 $Y=522220
X130 1237 66 1194 2 1 84 QDFFRBN $T=481740 527640 1 180 $X=469960 $Y=527260
X131 1219 66 1194 2 1 83 QDFFRBN $T=482360 537720 0 180 $X=470580 $Y=532300
X132 1249 61 1212 2 1 916 QDFFRBN $T=482980 507480 1 180 $X=471200 $Y=507100
X133 1250 61 70 2 1 1192 QDFFRBN $T=483600 396600 1 180 $X=471820 $Y=396220
X134 1213 61 1202 2 1 1251 QDFFRBN $T=472440 406680 0 0 $X=472440 $Y=406300
X135 1217 61 1202 2 1 1258 QDFFRBN $T=473060 426840 1 0 $X=473060 $Y=421420
X136 88 61 1212 2 1 784 QDFFRBN $T=492280 517560 0 180 $X=480500 $Y=512140
X137 1246 61 1267 2 1 1273 QDFFRBN $T=481120 426840 0 0 $X=481120 $Y=426460
X138 1275 61 1253 2 1 1024 QDFFRBN $T=492900 497400 1 180 $X=481120 $Y=497020
X139 1252 61 1267 2 1 1265 QDFFRBN $T=481740 436920 0 0 $X=481740 $Y=436540
X140 89 61 1253 2 1 810 QDFFRBN $T=494140 517560 1 180 $X=482360 $Y=517180
X141 1274 66 1194 2 1 87 QDFFRBN $T=494140 527640 1 180 $X=482360 $Y=527260
X142 90 61 1212 2 1 804 QDFFRBN $T=495380 507480 0 180 $X=483600 $Y=502060
X143 91 66 1194 2 1 809 QDFFRBN $T=495380 537720 0 180 $X=483600 $Y=532300
X144 1259 61 1202 2 1 1290 QDFFRBN $T=484840 406680 0 0 $X=484840 $Y=406300
X145 93 66 1253 2 1 972 QDFFRBN $T=497860 527640 0 180 $X=486080 $Y=522220
X146 1271 61 1293 2 1 1302 QDFFRBN $T=490420 457080 0 0 $X=490420 $Y=456700
X147 1278 61 1293 2 1 1299 QDFFRBN $T=492280 447000 0 0 $X=492280 $Y=446620
X148 96 61 1286 2 1 879 QDFFRBN $T=504060 477240 0 180 $X=492280 $Y=471820
X149 97 61 1287 2 1 998 QDFFRBN $T=504060 507480 1 180 $X=492280 $Y=507100
X150 1281 61 1298 2 1 1304 QDFFRBN $T=492900 436920 1 0 $X=492900 $Y=431500
X151 1307 61 1286 2 1 1276 QDFFRBN $T=504680 467160 0 180 $X=492900 $Y=461740
X152 103 61 1282 2 1 1009 QDFFRBN $T=507160 497400 0 180 $X=495380 $Y=491980
X153 109 61 1282 2 1 993 QDFFRBN $T=507160 497400 1 180 $X=495380 $Y=497020
X154 1288 66 1287 2 1 1319 QDFFRBN $T=495380 527640 0 0 $X=495380 $Y=527260
X155 1289 66 1287 2 1 1316 QDFFRBN $T=496000 517560 0 0 $X=496000 $Y=517180
X156 1270 61 1267 2 1 1325 QDFFRBN $T=499100 416760 1 0 $X=499100 $Y=411340
X157 1277 61 1267 2 1 1292 QDFFRBN $T=499100 416760 0 0 $X=499100 $Y=416380
X158 1291 61 1298 2 1 1321 QDFFRBN $T=499100 426840 0 0 $X=499100 $Y=426460
X159 1312 61 112 2 1 1338 QDFFRBN $T=506540 507480 0 0 $X=506540 $Y=507100
X160 1317 61 1335 2 1 1339 QDFFRBN $T=509020 477240 0 0 $X=509020 $Y=476860
X161 1318 61 1282 2 1 1341 QDFFRBN $T=509020 507480 1 0 $X=509020 $Y=502060
X162 1322 61 1335 2 1 1343 QDFFRBN $T=509640 467160 0 0 $X=509640 $Y=466780
X163 1323 61 1335 2 1 1344 QDFFRBN $T=509640 487320 0 0 $X=509640 $Y=486940
X164 1324 66 112 2 1 1347 QDFFRBN $T=509640 517560 0 0 $X=509640 $Y=517180
X165 1311 61 1293 2 1 1350 QDFFRBN $T=510260 447000 1 0 $X=510260 $Y=441580
X166 1326 61 1293 2 1 1348 QDFFRBN $T=510260 447000 0 0 $X=510260 $Y=446620
X167 1306 61 1293 2 1 1351 QDFFRBN $T=510880 457080 0 0 $X=510880 $Y=456700
X168 1354 66 116 2 1 1392 QDFFRBN $T=522660 517560 0 0 $X=522660 $Y=517180
X169 121 61 1386 2 1 1403 QDFFRBN $T=523900 497400 1 0 $X=523900 $Y=491980
X170 122 61 1386 2 1 1400 QDFFRBN $T=524520 487320 0 0 $X=524520 $Y=486940
X171 1365 61 1386 2 1 1406 QDFFRBN $T=525140 487320 1 0 $X=525140 $Y=481900
X172 1414 66 116 2 1 1380 QDFFRBN $T=542500 537720 0 180 $X=530720 $Y=532300
X173 1398 66 1417 2 1 1431 QDFFRBN $T=535060 527640 1 0 $X=535060 $Y=522220
X174 142 66 1417 2 1 1401 QDFFRBN $T=547460 517560 1 180 $X=535680 $Y=517180
X175 132 61 1386 2 1 1434 QDFFRBN $T=537540 487320 0 0 $X=537540 $Y=486940
X176 133 61 1386 2 1 1439 QDFFRBN $T=537540 497400 1 0 $X=537540 $Y=491980
X177 136 61 1386 2 1 1436 QDFFRBN $T=538780 497400 0 0 $X=538780 $Y=497020
X178 138 61 1377 2 1 1437 QDFFRBN $T=538780 507480 0 0 $X=538780 $Y=507100
X179 1422 61 1377 2 1 1444 QDFFRBN $T=539400 507480 1 0 $X=539400 $Y=502060
X180 1465 66 116 2 1 1426 QDFFRBN $T=554280 537720 0 180 $X=542500 $Y=532300
X181 146 66 1467 2 1 1408 QDFFRBN $T=549320 527640 1 0 $X=549320 $Y=522220
X182 147 66 1417 2 1 1438 QDFFRBN $T=549940 527640 0 0 $X=549940 $Y=527260
X183 1488 159 1467 2 1 1384 QDFFRBN $T=565440 517560 0 180 $X=553660 $Y=512140
X184 1499 159 1525 2 1 1545 QDFFRBN $T=561100 537720 1 0 $X=561100 $Y=532300
X185 169 159 1525 2 1 1385 QDFFRBN $T=574740 517560 1 180 $X=562960 $Y=517180
X186 1617 159 1525 2 1 1495 QDFFRBN $T=585280 527640 1 180 $X=573500 $Y=527260
X187 1555 159 173 2 1 1607 QDFFRBN $T=574120 537720 0 0 $X=574120 $Y=537340
X188 183 159 182 2 1 1623 QDFFRBN $T=617520 537720 1 180 $X=605740 $Y=537340
X189 185 159 1762 2 1 1780 QDFFRBN $T=618760 527640 0 0 $X=618760 $Y=527260
X190 190 159 187 2 1 1740 QDFFRBN $T=631160 537720 1 180 $X=619380 $Y=537340
X191 1796 159 1762 2 1 1422 QDFFRBN $T=637980 527640 0 180 $X=626200 $Y=522220
X192 1814 159 1762 2 1 1745 QDFFRBN $T=642320 537720 0 180 $X=630540 $Y=532300
X193 1824 159 1762 2 1 1617 QDFFRBN $T=644180 527640 1 180 $X=632400 $Y=527260
X194 1829 159 1762 2 1 1407 QDFFRBN $T=644800 517560 0 180 $X=633020 $Y=512140
X195 194 159 192 2 1 1843 QDFFRBN $T=636120 537720 0 0 $X=636120 $Y=537340
X196 202 204 215 2 1 220 QDFFRBN $T=648520 396600 1 0 $X=648520 $Y=391180
X197 203 204 215 2 1 224 QDFFRBN $T=649140 396600 0 0 $X=649140 $Y=396220
X198 207 204 215 2 1 222 QDFFRBN $T=651000 406680 1 0 $X=651000 $Y=401260
X199 208 204 215 2 1 1895 QDFFRBN $T=652240 406680 0 0 $X=652240 $Y=406300
X200 209 204 1885 2 1 1891 QDFFRBN $T=652860 426840 1 0 $X=652860 $Y=421420
X201 211 204 1885 2 1 1898 QDFFRBN $T=654100 426840 0 0 $X=654100 $Y=426460
X202 213 204 1888 2 1 1897 QDFFRBN $T=654720 477240 0 0 $X=654720 $Y=476860
X203 1876 204 1890 2 1 1901 QDFFRBN $T=655340 467160 0 0 $X=655340 $Y=466780
X204 216 204 1892 2 1 1899 QDFFRBN $T=655960 507480 1 0 $X=655960 $Y=502060
X205 1880 204 1888 2 1 1910 QDFFRBN $T=656580 487320 0 0 $X=656580 $Y=486940
X206 1863 204 1894 2 1 1883 QDFFRBN $T=656580 507480 0 0 $X=656580 $Y=507100
X207 1877 159 1894 2 1 1887 QDFFRBN $T=656580 517560 0 0 $X=656580 $Y=517180
X208 1878 159 1894 2 1 1903 QDFFRBN $T=656580 527640 1 0 $X=656580 $Y=522220
X209 217 204 1888 2 1 1952 QDFFRBN $T=657200 497400 1 0 $X=657200 $Y=491980
X210 1864 159 228 2 1 1881 QDFFRBN $T=657200 537720 0 0 $X=657200 $Y=537340
X211 1887 204 1896 2 1 1918 QDFFRBN $T=661540 457080 0 0 $X=661540 $Y=456700
X212 1912 159 1894 2 1 1687 QDFFRBN $T=673320 537720 0 180 $X=661540 $Y=532300
X213 225 204 1896 2 1 1927 QDFFRBN $T=663400 447000 0 0 $X=663400 $Y=446620
X214 226 204 1896 2 1 1915 QDFFRBN $T=664020 467160 1 0 $X=664020 $Y=461740
X215 227 204 1888 2 1 1932 QDFFRBN $T=664640 487320 1 0 $X=664640 $Y=481900
X216 1652 232 240 2 1 1946 QDFFRBN $T=666500 517560 1 0 $X=666500 $Y=512140
X217 1903 232 1890 2 1 1951 QDFFRBN $T=668980 507480 1 0 $X=668980 $Y=502060
X218 1831 232 1892 2 1 1963 QDFFRBN $T=669600 507480 0 0 $X=669600 $Y=507100
X219 1870 204 1890 2 1 1956 QDFFRBN $T=670220 487320 0 0 $X=670220 $Y=486940
X220 1766 159 240 2 1 1964 QDFFRBN $T=670220 517560 0 0 $X=670220 $Y=517180
X221 1917 159 1894 2 1 1935 QDFFRBN $T=670840 527640 0 0 $X=670840 $Y=527260
X222 1935 204 1890 2 1 1979 QDFFRBN $T=676420 497400 0 0 $X=676420 $Y=497020
X223 248 159 1987 2 1 2012 QDFFRBN $T=682620 537720 1 0 $X=682620 $Y=532300
X224 1871 232 1892 2 1 2024 QDFFRBN $T=683860 507480 0 0 $X=683860 $Y=507100
X225 1804 232 1892 2 1 2032 QDFFRBN $T=684480 517560 0 0 $X=684480 $Y=517180
X226 1685 159 1987 2 1 2036 QDFFRBN $T=684480 527640 0 0 $X=684480 $Y=527260
X227 253 232 1993 2 1 2029 QDFFRBN $T=686340 517560 1 0 $X=686340 $Y=512140
X228 1736 232 1987 2 1 2053 QDFFRBN $T=690060 527640 1 0 $X=690060 $Y=522220
X229 2030 232 1987 2 1 2098 QDFFRBN $T=696260 537720 1 0 $X=696260 $Y=532300
X230 2002 232 1993 2 1 2085 QDFFRBN $T=697500 507480 0 0 $X=697500 $Y=507100
X231 2045 232 1993 2 1 2100 QDFFRBN $T=698740 507480 1 0 $X=698740 $Y=502060
X232 262 232 1987 2 1 2086 QDFFRBN $T=698740 527640 0 0 $X=698740 $Y=527260
X233 263 232 1993 2 1 2112 QDFFRBN $T=699360 517560 1 0 $X=699360 $Y=512140
X234 266 232 1987 2 1 2120 QDFFRBN $T=701220 537720 0 0 $X=701220 $Y=537340
X235 2311 204 2332 2 1 2367 QDFFRBN $T=748960 497400 0 0 $X=748960 $Y=497020
X236 2340 204 2332 2 1 2315 QDFFRBN $T=762600 487320 1 180 $X=750820 $Y=486940
X237 2304 204 2332 2 1 2320 QDFFRBN $T=763220 497400 0 180 $X=751440 $Y=491980
X238 2394 204 2332 2 1 2351 QDFFRBN $T=769420 487320 0 180 $X=757640 $Y=481900
X239 2329 204 2332 2 1 2420 QDFFRBN $T=763220 497400 0 0 $X=763220 $Y=497020
X240 1874 204 2332 2 1 2453 QDFFRBN $T=769420 487320 1 0 $X=769420 $Y=481900
X241 1884 204 2444 2 1 2466 QDFFRBN $T=770660 467160 0 0 $X=770660 $Y=466780
X242 2407 204 2444 2 1 2489 QDFFRBN $T=770660 477240 1 0 $X=770660 $Y=471820
X243 2442 204 2479 2 1 2484 QDFFRBN $T=778100 497400 0 0 $X=778100 $Y=497020
X244 2446 204 2479 2 1 2493 QDFFRBN $T=778720 497400 1 0 $X=778720 $Y=491980
X245 2459 204 2469 2 1 2452 QDFFRBN $T=792360 467160 0 180 $X=780580 $Y=461740
X246 2488 204 2469 2 1 2457 QDFFRBN $T=792980 457080 0 180 $X=781200 $Y=451660
X247 2492 232 2479 2 1 2462 QDFFRBN $T=794220 507480 0 180 $X=782440 $Y=502060
X248 1813 204 2469 2 1 2533 QDFFRBN $T=791120 436920 1 0 $X=791120 $Y=431500
X249 2464 204 2510 2 1 2513 QDFFRBN $T=791740 416760 1 0 $X=791740 $Y=411340
X250 2501 204 2469 2 1 2538 QDFFRBN $T=792360 447000 0 0 $X=792360 $Y=446620
X251 2507 232 2479 2 1 2532 QDFFRBN $T=792980 497400 0 0 $X=792980 $Y=497020
X252 2188 232 322 2 1 329 QDFFRBN $T=794220 527640 1 0 $X=794220 $Y=522220
X253 2225 232 322 2 1 328 QDFFRBN $T=794220 537720 1 0 $X=794220 $Y=532300
X254 331 232 2520 2 1 2514 QDFFRBN $T=808480 507480 1 180 $X=796700 $Y=507100
X255 2388 232 2560 2 1 339 QDFFRBN $T=802900 527640 0 0 $X=802900 $Y=527260
X256 773 232 337 2 1 2593 QDFFRBN $T=806000 537720 1 0 $X=806000 $Y=532300
X257 2374 232 337 2 1 341 QDFFRBN $T=808480 537720 0 0 $X=808480 $Y=537340
X258 343 232 2576 2 1 2555 QDFFRBN $T=821500 497400 0 180 $X=809720 $Y=491980
X259 2447 232 2560 2 1 348 QDFFRBN $T=813440 517560 0 0 $X=813440 $Y=517180
X260 875 232 2560 2 1 2634 QDFFRBN $T=813440 527640 1 0 $X=813440 $Y=522220
X261 2642 344 340 2 1 338 QDFFRBN $T=827080 396600 0 180 $X=815300 $Y=391180
X262 696 232 346 2 1 2653 QDFFRBN $T=817780 537720 1 0 $X=817780 $Y=532300
X263 610 232 346 2 1 2671 QDFFRBN $T=822120 537720 0 0 $X=822120 $Y=537340
X264 2624 232 2670 2 1 2687 QDFFRBN $T=825220 487320 0 0 $X=825220 $Y=486940
X265 2546 232 2670 2 1 2681 QDFFRBN $T=825220 497400 1 0 $X=825220 $Y=491980
X266 871 232 2670 2 1 2689 QDFFRBN $T=825220 497400 0 0 $X=825220 $Y=497020
X267 347 232 2670 2 1 2705 QDFFRBN $T=825840 507480 1 0 $X=825840 $Y=502060
X268 2509 232 2670 2 1 2682 QDFFRBN $T=827080 507480 0 0 $X=827080 $Y=507100
X269 352 344 340 2 1 2642 QDFFRBN $T=839480 396600 0 180 $X=827700 $Y=391180
X270 2494 232 2670 2 1 353 QDFFRBN $T=827700 517560 1 0 $X=827700 $Y=512140
X271 2472 232 2679 2 1 354 QDFFRBN $T=827700 527640 1 0 $X=827700 $Y=522220
X272 2649 344 2706 2 1 2730 QDFFRBN $T=834520 487320 1 0 $X=834520 $Y=481900
X273 2608 344 2706 2 1 2722 QDFFRBN $T=835760 477240 0 0 $X=835760 $Y=476860
X274 2697 344 2712 2 1 367 QDFFRBN $T=840720 467160 1 0 $X=840720 $Y=461740
X275 2680 344 2706 2 1 366 QDFFRBN $T=840720 477240 1 0 $X=840720 $Y=471820
X276 2711 344 2731 2 1 2749 QDFFRBN $T=843200 416760 1 0 $X=843200 $Y=411340
X277 2757 344 358 2 1 363 QDFFRBN $T=858700 396600 0 180 $X=846920 $Y=391180
X278 2672 344 2706 2 1 369 QDFFRBN $T=847540 477240 0 0 $X=847540 $Y=476860
X279 2740 344 2731 2 1 2711 QDFFRBN $T=859940 426840 0 180 $X=848160 $Y=421420
X280 2737 344 2754 2 1 2769 QDFFRBN $T=853120 447000 1 0 $X=853120 $Y=441580
X281 2769 344 2712 2 1 2734 QDFFRBN $T=864900 457080 0 180 $X=853120 $Y=451660
X282 2772 344 2717 2 1 2740 QDFFRBN $T=865520 426840 1 180 $X=853740 $Y=426460
X283 2743 344 2717 2 1 2772 QDFFRBN $T=854360 436920 1 0 $X=854360 $Y=431500
X284 2777 344 2754 2 1 2737 QDFFRBN $T=866760 447000 1 180 $X=854980 $Y=446620
X285 2746 344 372 2 1 2709 QDFFRBN $T=855600 406680 1 0 $X=855600 $Y=401260
X286 2611 344 2754 2 1 377 QDFFRBN $T=856220 467160 1 0 $X=856220 $Y=461740
X287 2683 344 2706 2 1 2828 QDFFRBN $T=857460 477240 1 0 $X=857460 $Y=471820
X288 2692 344 2706 2 1 380 QDFFRBN $T=859320 477240 0 0 $X=859320 $Y=476860
X289 2804 344 372 2 1 2757 QDFFRBN $T=872960 396600 0 180 $X=861180 $Y=391180
X290 2783 344 2770 2 1 2791 QDFFRBN $T=866140 416760 0 0 $X=866140 $Y=416380
X291 2695 344 2784 2 1 2823 QDFFRBN $T=866760 447000 1 0 $X=866760 $Y=441580
X292 2789 2813 2770 2 1 2783 QDFFRBN $T=879160 426840 0 180 $X=867380 $Y=421420
X293 2819 344 2797 2 1 2777 QDFFRBN $T=879780 457080 0 180 $X=868000 $Y=451660
X294 2791 344 2770 2 1 2822 QDFFRBN $T=868620 416760 1 0 $X=868620 $Y=411340
X295 2851 2813 2784 2 1 2789 QDFFRBN $T=880400 436920 0 180 $X=868620 $Y=431500
X296 2832 2813 2784 2 1 2790 QDFFRBN $T=880400 436920 1 180 $X=868620 $Y=436540
X297 2790 344 2797 2 1 2819 QDFFRBN $T=868620 447000 0 0 $X=868620 $Y=446620
X298 2721 344 2797 2 1 388 QDFFRBN $T=868620 457080 0 0 $X=868620 $Y=456700
X299 2710 344 2797 2 1 394 QDFFRBN $T=869240 467160 1 0 $X=869240 $Y=461740
X300 2678 344 2785 2 1 2837 QDFFRBN $T=869860 467160 0 0 $X=869860 $Y=466780
X301 2696 344 2785 2 1 390 QDFFRBN $T=871100 477240 0 0 $X=871100 $Y=476860
X302 2836 391 372 2 1 2804 QDFFRBN $T=885980 396600 0 180 $X=874200 $Y=391180
X303 2847 2813 2770 2 1 383 QDFFRBN $T=889700 406680 1 180 $X=877920 $Y=406300
X304 2833 2813 2797 2 1 2880 QDFFRBN $T=881020 447000 1 0 $X=881020 $Y=441580
X305 2829 2813 2785 2 1 2830 QDFFRBN $T=892800 457080 0 180 $X=881020 $Y=451660
X306 2880 2813 2797 2 1 2832 QDFFRBN $T=893420 436920 1 180 $X=881640 $Y=436540
X307 2830 2813 2785 2 1 2897 QDFFRBN $T=882260 457080 0 0 $X=882260 $Y=456700
X308 2886 2813 395 2 1 2840 QDFFRBN $T=894660 406680 0 180 $X=882880 $Y=401260
X309 2843 2813 2877 2 1 2898 QDFFRBN $T=882880 467160 0 0 $X=882880 $Y=466780
X310 2844 2813 2877 2 1 2889 QDFFRBN $T=882880 477240 0 0 $X=882880 $Y=476860
X311 2840 391 395 2 1 2925 QDFFRBN $T=883500 396600 0 0 $X=883500 $Y=396220
X312 2903 2813 395 2 1 2847 QDFFRBN $T=895280 416760 0 180 $X=883500 $Y=411340
X313 2917 2813 2890 2 1 2851 QDFFRBN $T=903340 436920 0 180 $X=891560 $Y=431500
X314 2883 2813 2909 2 1 2928 QDFFRBN $T=892180 487320 1 0 $X=892180 $Y=481900
X315 2925 391 395 2 1 402 QDFFRBN $T=905200 396600 0 180 $X=893420 $Y=391180
X316 2930 391 395 2 1 2886 QDFFRBN $T=906440 406680 0 180 $X=894660 $Y=401260
X317 2889 2813 2900 2 1 2883 QDFFRBN $T=894660 477240 0 0 $X=894660 $Y=476860
X318 2897 2813 2900 2 1 2941 QDFFRBN $T=895900 457080 0 0 $X=895900 $Y=456700
X319 2898 2813 2900 2 1 2952 QDFFRBN $T=895900 467160 0 0 $X=895900 $Y=466780
X320 2941 2813 2890 2 1 2902 QDFFRBN $T=909540 457080 0 180 $X=897760 $Y=451660
X321 2928 2813 2909 2 1 2963 QDFFRBN $T=903960 487320 1 0 $X=903960 $Y=481900
X322 2959 2813 2890 2 1 2903 QDFFRBN $T=916360 436920 0 180 $X=904580 $Y=431500
X323 418 391 2922 2 1 2929 QDFFRBN $T=917600 406680 1 180 $X=905820 $Y=406300
X324 2973 2813 2950 2 1 2934 QDFFRBN $T=918840 447000 0 180 $X=907060 $Y=441580
X325 2940 391 417 2 1 423 QDFFRBN $T=907680 396600 1 0 $X=907680 $Y=391180
X326 2914 2813 2950 2 1 3015 QDFFRBN $T=907680 447000 0 0 $X=907680 $Y=446620
X327 2998 2813 2950 2 1 2959 QDFFRBN $T=923800 436920 1 180 $X=912020 $Y=436540
X328 2966 2813 2909 2 1 2997 QDFFRBN $T=912020 457080 0 0 $X=912020 $Y=456700
X329 3020 2813 2986 2 1 2966 QDFFRBN $T=925660 457080 0 180 $X=913880 $Y=451660
X330 3040 2813 2909 2 1 2978 QDFFRBN $T=928140 487320 0 180 $X=916360 $Y=481900
X331 3033 2813 3003 2 1 2985 QDFFRBN $T=928760 426840 0 180 $X=916980 $Y=421420
X332 2952 2813 2909 2 1 3040 QDFFRBN $T=918220 477240 0 0 $X=918220 $Y=476860
X333 3007 391 417 2 1 2940 QDFFRBN $T=932480 396600 0 180 $X=920700 $Y=391180
X334 3058 391 2922 2 1 3007 QDFFRBN $T=933100 396600 1 180 $X=921320 $Y=396220
X335 2971 2813 3034 2 1 3033 QDFFRBN $T=921320 436920 1 0 $X=921320 $Y=431500
X336 3066 2813 3003 2 1 3024 QDFFRBN $T=936820 416760 0 180 $X=925040 $Y=411340
X337 3061 2813 3034 2 1 2971 QDFFRBN $T=937440 436920 1 180 $X=925660 $Y=436540
X338 3015 2813 3051 2 1 3020 QDFFRBN $T=925660 457080 1 0 $X=925660 $Y=451660
X339 3022 2813 3034 2 1 3061 QDFFRBN $T=926900 447000 1 0 $X=926900 $Y=441580
X340 2985 2813 3003 2 1 3066 QDFFRBN $T=928760 426840 1 0 $X=928760 $Y=421420
X341 2984 2813 3052 2 1 3056 QDFFRBN $T=930000 497400 1 0 $X=930000 $Y=491980
X342 3050 2813 3052 2 1 3076 QDFFRBN $T=931240 487320 0 0 $X=931240 $Y=486940
X343 3047 2813 3052 2 1 3059 QDFFRBN $T=931240 507480 1 0 $X=931240 $Y=502060
X344 3073 2813 3051 2 1 3048 QDFFRBN $T=943640 467160 0 180 $X=931860 $Y=461740
X345 3076 2813 3051 2 1 3049 QDFFRBN $T=943640 477240 0 180 $X=931860 $Y=471820
X346 3048 2813 3051 2 1 3080 QDFFRBN $T=934340 457080 0 0 $X=934340 $Y=456700
X347 3056 2813 3052 2 1 3086 QDFFRBN $T=934340 477240 0 0 $X=934340 $Y=476860
X348 3059 2813 3052 2 1 3073 QDFFRBN $T=935580 487320 1 0 $X=935580 $Y=481900
X349 433 2813 431 2 1 3060 QDFFRBN $T=947980 527640 1 180 $X=936200 $Y=527260
X350 3060 430 431 2 1 3087 QDFFRBN $T=936820 537720 1 0 $X=936820 $Y=532300
X351 3062 2813 3079 2 1 3084 QDFFRBN $T=937440 447000 0 0 $X=937440 $Y=446620
X352 3049 2813 3051 2 1 3062 QDFFRBN $T=949840 457080 0 180 $X=938060 $Y=451660
X353 3064 2813 3081 2 1 3099 QDFFRBN $T=938060 527640 1 0 $X=938060 $Y=522220
X354 3065 2813 3081 2 1 3106 QDFFRBN $T=938680 517560 0 0 $X=938680 $Y=517180
X355 3098 2813 3052 2 1 3068 QDFFRBN $T=951700 497400 1 180 $X=939920 $Y=497020
X356 3083 2813 3079 2 1 3070 QDFFRBN $T=952320 436920 1 180 $X=940540 $Y=436540
X357 2904 2813 3081 2 1 3071 QDFFRBN $T=952320 517560 0 180 $X=940540 $Y=512140
X358 3071 2813 3081 2 1 3098 QDFFRBN $T=941160 507480 0 0 $X=941160 $Y=507100
X359 3108 391 3075 2 1 3077 QDFFRBN $T=954180 406680 0 180 $X=942400 $Y=401260
X360 3074 2813 3075 2 1 3108 QDFFRBN $T=943020 406680 0 0 $X=943020 $Y=406300
X361 3068 2813 2953 2 1 3110 QDFFRBN $T=943020 497400 1 0 $X=943020 $Y=491980
X362 3082 2813 3079 2 1 3118 QDFFRBN $T=943640 447000 1 0 $X=943640 $Y=441580
X363 3118 2813 3079 2 1 3083 QDFFRBN $T=957280 436920 0 180 $X=945500 $Y=431500
X364 3099 2813 3081 2 1 3065 QDFFRBN $T=951700 517560 0 0 $X=951700 $Y=517180
X365 3106 2813 3081 2 1 3150 QDFFRBN $T=951700 527640 1 0 $X=951700 $Y=522220
X366 3167 3151 3134 2 1 3112 QDFFRBN $T=967200 426840 1 180 $X=955420 $Y=426460
X367 3114 2813 3134 2 1 3167 QDFFRBN $T=955420 436920 0 0 $X=955420 $Y=436540
X368 3124 391 3164 2 1 3180 QDFFRBN $T=957280 396600 0 0 $X=957280 $Y=396220
X369 3091 2813 3163 2 1 3186 QDFFRBN $T=957900 447000 1 0 $X=957900 $Y=441580
X370 3180 391 440 2 1 442 QDFFRBN $T=970920 396600 0 180 $X=959140 $Y=391180
X371 3145 3151 3173 2 1 3188 QDFFRBN $T=959760 457080 0 0 $X=959760 $Y=456700
X372 3179 3151 2953 2 1 3149 QDFFRBN $T=972780 487320 0 180 $X=961000 $Y=481900
X373 3152 3151 2953 2 1 3189 QDFFRBN $T=961000 497400 1 0 $X=961000 $Y=491980
X374 3149 3151 2953 2 1 3152 QDFFRBN $T=973400 487320 1 180 $X=961620 $Y=486940
X375 3157 430 3169 2 1 3196 QDFFRBN $T=965340 517560 0 0 $X=965340 $Y=517180
X376 3158 430 3169 2 1 3195 QDFFRBN $T=965340 527640 1 0 $X=965340 $Y=522220
X377 3175 3151 3163 2 1 3197 QDFFRBN $T=967820 436920 1 0 $X=967820 $Y=431500
X378 3197 3151 3163 2 1 3177 QDFFRBN $T=980840 426840 1 180 $X=969060 $Y=426460
X379 3205 3151 3163 2 1 3175 QDFFRBN $T=980840 436920 1 180 $X=969060 $Y=436540
X380 449 3151 3171 2 1 3179 QDFFRBN $T=980840 477240 1 180 $X=969060 $Y=476860
X381 3182 391 3161 2 1 3198 QDFFRBN $T=969680 406680 1 0 $X=969680 $Y=401260
X382 3148 3151 3171 2 1 3203 QDFFRBN $T=969680 477240 1 0 $X=969680 $Y=471820
X383 3198 446 3164 2 1 3184 QDFFRBN $T=982080 396600 1 180 $X=970300 $Y=396220
X384 3181 3151 3192 2 1 3205 QDFFRBN $T=970920 447000 0 0 $X=970920 $Y=446620
X385 3203 3151 3171 2 1 3165 QDFFRBN $T=982700 467160 1 180 $X=970920 $Y=466780
X386 3207 3151 3192 2 1 3145 QDFFRBN $T=983320 457080 0 180 $X=971540 $Y=451660
X387 3188 3151 3173 2 1 3162 QDFFRBN $T=983320 457080 1 180 $X=971540 $Y=456700
X388 447 3151 3194 2 1 3209 QDFFRBN $T=971540 507480 0 0 $X=971540 $Y=507100
X389 3125 3151 3194 2 1 3216 QDFFRBN $T=971540 517560 1 0 $X=971540 $Y=512140
X390 3184 391 450 2 1 452 QDFFRBN $T=972160 396600 1 0 $X=972160 $Y=391180
X391 3209 3151 3194 2 1 3191 QDFFRBN $T=985180 507480 0 180 $X=973400 $Y=502060
X392 3174 430 451 2 1 3219 QDFFRBN $T=975260 537720 1 0 $X=975260 $Y=532300
X393 454 430 451 2 1 448 QDFFRBN $T=988900 537720 1 180 $X=977120 $Y=537340
X394 3196 430 3169 2 1 3187 QDFFRBN $T=989520 527640 0 180 $X=977740 $Y=522220
X395 3191 3151 3211 2 1 3225 QDFFRBN $T=978360 487320 0 0 $X=978360 $Y=486940
X396 3202 3151 3211 2 1 3230 QDFFRBN $T=980220 487320 1 0 $X=980220 $Y=481900
X397 3225 3151 3211 2 1 3193 QDFFRBN $T=993240 497400 0 180 $X=981460 $Y=491980
X398 3195 3151 3194 2 1 3215 QDFFRBN $T=981460 517560 0 0 $X=981460 $Y=517180
X399 3186 3151 3192 2 1 3214 QDFFRBN $T=982700 436920 0 0 $X=982700 $Y=436540
X400 457 446 3204 2 1 3206 QDFFRBN $T=995100 406680 0 180 $X=983320 $Y=401260
X401 3208 3151 3192 2 1 3231 QDFFRBN $T=983320 447000 1 0 $X=983320 $Y=441580
X402 3228 3151 3171 2 1 3148 QDFFRBN $T=995100 477240 0 180 $X=983320 $Y=471820
X403 2943 3151 3173 2 1 3207 QDFFRBN $T=995720 457080 0 180 $X=983940 $Y=451660
X404 3178 3151 3173 2 1 3208 QDFFRBN $T=995720 457080 1 180 $X=983940 $Y=456700
X405 3214 446 3204 2 1 3233 QDFFRBN $T=985180 416760 1 0 $X=985180 $Y=411340
X406 3215 3151 3194 2 1 3247 QDFFRBN $T=985180 507480 0 0 $X=985180 $Y=507100
X407 3216 3151 3194 2 1 3236 QDFFRBN $T=985180 517560 1 0 $X=985180 $Y=512140
X408 3219 430 451 2 1 3239 QDFFRBN $T=987040 537720 1 0 $X=987040 $Y=532300
X409 3200 3151 3224 2 1 3254 QDFFRBN $T=990760 487320 0 0 $X=990760 $Y=486940
X410 2891 3151 3224 2 1 3228 QDFFRBN $T=1003780 477240 1 180 $X=992000 $Y=476860
X411 3230 3151 3224 2 1 3249 QDFFRBN $T=993860 487320 1 0 $X=993860 $Y=481900
X412 3231 446 3252 2 1 3235 QDFFRBN $T=994480 426840 1 0 $X=994480 $Y=421420
X413 3249 3151 3238 2 1 3232 QDFFRBN $T=1006880 467160 0 180 $X=995100 $Y=461740
X414 3235 446 3252 2 1 3264 QDFFRBN $T=995720 416760 0 0 $X=995720 $Y=416380
X415 3232 3151 3238 2 1 3268 QDFFRBN $T=996960 457080 0 0 $X=996960 $Y=456700
X416 3240 446 450 2 1 471 QDFFRBN $T=997580 396600 0 0 $X=997580 $Y=396220
X417 3272 3151 3250 2 1 3244 QDFFRBN $T=1010600 497400 1 180 $X=998820 $Y=497020
X418 3244 3151 3250 2 1 3273 QDFFRBN $T=1000680 497400 1 0 $X=1000680 $Y=491980
X419 3254 3151 3224 2 1 3265 QDFFRBN $T=1003780 487320 0 0 $X=1003780 $Y=486940
X420 3279 3151 3252 2 1 3256 QDFFRBN $T=1018660 426840 0 180 $X=1006880 $Y=421420
X421 3281 3151 3238 2 1 3258 QDFFRBN $T=1018660 457080 0 180 $X=1006880 $Y=451660
X422 3287 430 472 2 1 469 QDFFRBN $T=1018660 537720 1 180 $X=1006880 $Y=537340
X423 3283 446 473 2 1 470 QDFFRBN $T=1019280 396600 0 180 $X=1007500 $Y=391180
X424 3259 446 3204 2 1 3283 QDFFRBN $T=1007500 406680 1 0 $X=1007500 $Y=401260
X425 3257 3151 3267 2 1 3279 QDFFRBN $T=1007500 436920 1 0 $X=1007500 $Y=431500
X426 3239 430 472 2 1 3285 QDFFRBN $T=1008120 527640 1 0 $X=1008120 $Y=522220
X427 3268 3151 3238 2 1 3281 QDFFRBN $T=1009360 457080 0 0 $X=1009360 $Y=456700
X428 3273 3151 3291 2 1 3300 QDFFRBN $T=1013080 497400 0 0 $X=1013080 $Y=497020
X429 3236 3151 3292 2 1 3274 QDFFRBN $T=1013080 517560 1 0 $X=1013080 $Y=512140
X430 3274 3151 3292 2 1 3299 QDFFRBN $T=1013700 507480 0 0 $X=1013700 $Y=507100
X431 3265 3151 3291 2 1 3282 QDFFRBN $T=1015560 497400 1 0 $X=1015560 $Y=491980
X432 3282 3151 3291 2 1 3301 QDFFRBN $T=1016800 487320 0 0 $X=1016800 $Y=486940
X433 3256 3151 3276 2 1 3295 QDFFRBN $T=1018660 426840 1 0 $X=1018660 $Y=421420
X434 3302 3151 3294 2 1 3286 QDFFRBN $T=1030440 467160 1 180 $X=1018660 $Y=466780
X435 3317 3151 3294 2 1 3277 QDFFRBN $T=1030440 477240 0 180 $X=1018660 $Y=471820
X436 3264 446 3276 2 1 3306 QDFFRBN $T=1019900 416760 1 0 $X=1019900 $Y=411340
X437 3286 3151 3294 2 1 3303 QDFFRBN $T=1019900 467160 1 0 $X=1019900 $Y=461740
X438 3305 3151 3267 2 1 3269 QDFFRBN $T=1032300 436920 1 180 $X=1020520 $Y=436540
X439 3289 446 475 2 1 477 QDFFRBN $T=1021140 396600 1 0 $X=1021140 $Y=391180
X440 3306 446 475 2 1 3289 QDFFRBN $T=1032920 406680 0 180 $X=1021140 $Y=401260
X441 479 446 3276 2 1 3260 QDFFRBN $T=1032920 406680 1 180 $X=1021140 $Y=406300
X442 3295 3151 3276 2 1 3310 QDFFRBN $T=1021760 426840 0 0 $X=1021760 $Y=426460
X443 3309 3151 3297 2 1 3278 QDFFRBN $T=1034160 517560 1 180 $X=1022380 $Y=517180
X444 3316 430 3297 2 1 3296 QDFFRBN $T=1034160 527640 0 180 $X=1022380 $Y=522220
X445 3300 3151 3291 2 1 3326 QDFFRBN $T=1026100 497400 0 0 $X=1026100 $Y=497020
X446 3299 3151 3297 2 1 3320 QDFFRBN $T=1026100 517560 1 0 $X=1026100 $Y=512140
X447 3304 3151 3315 2 1 3333 QDFFRBN $T=1030440 416760 0 0 $X=1030440 $Y=416380
X448 3329 3151 3315 2 1 3304 QDFFRBN $T=1042840 426840 0 180 $X=1031060 $Y=421420
X449 3308 446 475 2 1 3328 QDFFRBN $T=1032300 396600 0 0 $X=1032300 $Y=396220
X450 3307 3151 481 2 1 3334 QDFFRBN $T=1032300 457080 0 0 $X=1032300 $Y=456700
X451 3310 3151 3315 2 1 3329 QDFFRBN $T=1033540 426840 0 0 $X=1033540 $Y=426460
X452 3313 3327 481 2 1 3312 QDFFRBN $T=1045320 447000 1 180 $X=1033540 $Y=446620
X453 3334 3327 481 2 1 3313 QDFFRBN $T=1045320 457080 0 180 $X=1033540 $Y=451660
X454 3338 446 475 2 1 3308 QDFFRBN $T=1045940 396600 0 180 $X=1034160 $Y=391180
X455 3312 3151 3330 2 1 3343 QDFFRBN $T=1034160 447000 1 0 $X=1034160 $Y=441580
X456 3337 430 3297 2 1 3316 QDFFRBN $T=1047180 527640 0 180 $X=1035400 $Y=522220
X457 3319 3151 3297 2 1 3337 QDFFRBN $T=1036020 517560 0 0 $X=1036020 $Y=517180
X458 3324 3327 3311 2 1 3346 QDFFRBN $T=1038500 487320 0 0 $X=1038500 $Y=486940
X459 484 430 482 2 1 3323 QDFFRBN $T=1051520 537720 1 180 $X=1039740 $Y=537340
X460 3323 430 476 2 1 3359 QDFFRBN $T=1040360 537720 1 0 $X=1040360 $Y=532300
X461 3331 3327 3330 2 1 3360 QDFFRBN $T=1042840 436920 1 0 $X=1042840 $Y=431500
X462 3366 3327 481 2 1 3332 QDFFRBN $T=1055860 467160 0 180 $X=1044080 $Y=461740
X463 3369 485 3336 2 1 3338 QDFFRBN $T=1058960 396600 0 180 $X=1047180 $Y=391180
X464 3352 486 3335 2 1 3370 QDFFRBN $T=1051520 517560 0 0 $X=1051520 $Y=517180
X465 3387 3327 3335 2 1 3352 QDFFRBN $T=1064540 517560 0 180 $X=1052760 $Y=512140
X466 3356 485 3364 2 1 3365 QDFFRBN $T=1053380 406680 0 0 $X=1053380 $Y=406300
X467 3357 3327 3371 2 1 3377 QDFFRBN $T=1053380 497400 0 0 $X=1053380 $Y=497020
X468 3376 486 482 2 1 487 QDFFRBN $T=1065160 537720 1 180 $X=1053380 $Y=537340
X469 3362 485 3364 2 1 3356 QDFFRBN $T=1065780 416760 0 180 $X=1054000 $Y=411340
X470 3359 486 482 2 1 3376 QDFFRBN $T=1054000 537720 1 0 $X=1054000 $Y=532300
X471 3379 3327 3335 2 1 3353 QDFFRBN $T=1066400 507480 1 180 $X=1054620 $Y=507100
X472 3383 3327 3368 2 1 3363 QDFFRBN $T=1068260 467160 1 180 $X=1056480 $Y=466780
X473 3363 3327 3368 2 1 3391 QDFFRBN $T=1057100 467160 1 0 $X=1057100 $Y=461740
X474 3380 3327 3350 2 1 3366 QDFFRBN $T=1073220 457080 0 180 $X=1061440 $Y=451660
X475 3374 3327 3371 2 1 3390 QDFFRBN $T=1061440 497400 1 0 $X=1061440 $Y=491980
X476 3392 3327 3371 2 1 3374 QDFFRBN $T=1073840 487320 0 180 $X=1062060 $Y=481900
X477 3375 3327 3368 2 1 3392 QDFFRBN $T=1062680 477240 0 0 $X=1062680 $Y=476860
X478 3373 486 3335 2 1 3404 QDFFRBN $T=1064540 517560 0 0 $X=1064540 $Y=517180
X479 3411 3327 3350 2 1 3380 QDFFRBN $T=1076940 447000 1 180 $X=1065160 $Y=446620
X480 3377 3327 3371 2 1 3426 QDFFRBN $T=1065160 507480 1 0 $X=1065160 $Y=502060
X481 3397 486 3386 2 1 3373 QDFFRBN $T=1076940 527640 0 180 $X=1065160 $Y=522220
X482 3398 3327 3371 2 1 3379 QDFFRBN $T=1077560 497400 1 180 $X=1065780 $Y=497020
X483 3384 486 3396 2 1 3397 QDFFRBN $T=1067020 527640 0 0 $X=1067020 $Y=527260
X484 3407 485 3364 2 1 3385 QDFFRBN $T=1079420 406680 1 180 $X=1067640 $Y=406300
X485 491 486 482 2 1 3384 QDFFRBN $T=1079420 537720 1 180 $X=1067640 $Y=537340
X486 3385 485 3393 2 1 3389 QDFFRBN $T=1068260 416760 1 0 $X=1068260 $Y=411340
X487 3389 485 3393 2 1 3410 QDFFRBN $T=1069500 426840 1 0 $X=1069500 $Y=421420
X488 3390 3327 3402 2 1 3400 QDFFRBN $T=1069500 487320 0 0 $X=1069500 $Y=486940
X489 3405 486 3386 2 1 3387 QDFFRBN $T=1081280 517560 0 180 $X=1069500 $Y=512140
X490 3423 3327 3395 2 1 3399 QDFFRBN $T=1088100 477240 0 180 $X=1076320 $Y=471820
X491 3400 3327 3395 2 1 3423 QDFFRBN $T=1076320 487320 1 0 $X=1076320 $Y=481900
X492 3399 3327 3395 2 1 3424 QDFFRBN $T=1076940 477240 0 0 $X=1076940 $Y=476860
X493 3429 3327 3402 2 1 3398 QDFFRBN $T=1088720 507480 1 180 $X=1076940 $Y=507100
X494 3404 486 3386 2 1 3425 QDFFRBN $T=1076940 517560 0 0 $X=1076940 $Y=517180
X495 3424 3327 3402 2 1 3403 QDFFRBN $T=1089340 497400 0 180 $X=1077560 $Y=491980
X496 3403 3327 3402 2 1 3357 QDFFRBN $T=1089340 497400 1 180 $X=1077560 $Y=497020
X497 3394 485 3417 2 1 3406 QDFFRBN $T=1079420 396600 1 0 $X=1079420 $Y=391180
X498 3406 485 3417 2 1 3436 QDFFRBN $T=1079420 396600 0 0 $X=1079420 $Y=396220
X499 3433 486 3386 2 1 3405 QDFFRBN $T=1091200 527640 0 180 $X=1079420 $Y=522220
X500 3409 486 3396 2 1 3433 QDFFRBN $T=1080040 537720 1 0 $X=1080040 $Y=532300
X501 493 486 492 2 1 3409 QDFFRBN $T=1093680 537720 1 180 $X=1081900 $Y=537340
X502 3414 3327 3428 2 1 3434 QDFFRBN $T=1082520 447000 0 0 $X=1082520 $Y=446620
X503 3420 485 3419 2 1 3438 QDFFRBN $T=1084380 426840 1 0 $X=1084380 $Y=421420
X504 3438 485 3417 2 1 3421 QDFFRBN $T=1097400 416760 1 180 $X=1085620 $Y=416380
X505 3427 486 3396 2 1 497 QDFFRBN $T=1088720 527640 0 0 $X=1088720 $Y=527260
X506 3421 485 3419 2 1 3451 QDFFRBN $T=1089340 416760 1 0 $X=1089340 $Y=411340
X507 3425 486 3386 2 1 3427 QDFFRBN $T=1101740 517560 1 180 $X=1089960 $Y=517180
X508 3447 3327 3402 2 1 3429 QDFFRBN $T=1102980 507480 1 180 $X=1091200 $Y=507100
X509 3432 3327 3431 2 1 3447 QDFFRBN $T=1091820 497400 0 0 $X=1091820 $Y=497020
X510 3461 3327 3431 2 1 3432 QDFFRBN $T=1104840 497400 0 180 $X=1093060 $Y=491980
X511 3453 485 3440 2 1 494 QDFFRBN $T=1106080 396600 0 180 $X=1094300 $Y=391180
X512 3456 486 496 2 1 495 QDFFRBN $T=1107940 537720 1 180 $X=1096160 $Y=537340
X513 3441 3327 3446 2 1 3458 QDFFRBN $T=1097400 447000 0 0 $X=1097400 $Y=446620
X514 3459 3327 3422 2 1 3443 QDFFRBN $T=1109180 467160 1 180 $X=1097400 $Y=466780
X515 3445 3327 3431 2 1 3461 QDFFRBN $T=1098020 487320 1 0 $X=1098020 $Y=481900
X516 3426 3327 3431 2 1 3465 QDFFRBN $T=1098020 507480 1 0 $X=1098020 $Y=502060
X517 3472 486 3386 2 1 3449 QDFFRBN $T=1113520 527640 0 180 $X=1101740 $Y=522220
X518 3465 3327 3455 2 1 3485 QDFFRBN $T=1111660 507480 1 0 $X=1111660 $Y=502060
X519 3463 3327 3446 2 1 3462 QDFFRBN $T=1124060 457080 0 180 $X=1112280 $Y=451660
X520 3482 3327 3476 2 1 3464 QDFFRBN $T=1124060 487320 0 180 $X=1112280 $Y=481900
X521 3469 3327 3476 2 1 3482 QDFFRBN $T=1112280 497400 1 0 $X=1112280 $Y=491980
X522 3470 485 3466 2 1 3471 QDFFRBN $T=1125300 416760 1 180 $X=1113520 $Y=416380
X523 3489 485 3466 2 1 3473 QDFFRBN $T=1125920 416760 0 180 $X=1114140 $Y=411340
X524 3471 485 3467 2 1 3484 QDFFRBN $T=1114140 426840 1 0 $X=1114140 $Y=421420
X525 3474 3327 3467 2 1 3475 QDFFRBN $T=1114140 436920 0 0 $X=1114140 $Y=436540
X526 3485 486 3476 2 1 3469 QDFFRBN $T=1127780 497400 1 180 $X=1116000 $Y=497020
X527 3486 486 3455 2 1 3477 QDFFRBN $T=1128400 517560 0 180 $X=1116620 $Y=512140
X528 499 486 498 2 1 3488 QDFFRBN $T=1116620 537720 0 0 $X=1116620 $Y=537340
X529 513 2 515 1 INV1S $T=303800 537720 1 0 $X=303800 $Y=532300
X530 523 2 518 1 INV1S $T=310620 507480 0 180 $X=309380 $Y=502060
X531 516 2 17 1 INV1S $T=310620 537720 0 0 $X=310620 $Y=537340
X532 536 2 529 1 INV1S $T=314340 487320 0 180 $X=313100 $Y=481900
X533 547 2 541 1 INV1S $T=319920 487320 0 180 $X=318680 $Y=481900
X534 546 2 549 1 INV1S $T=319300 477240 0 0 $X=319300 $Y=476860
X535 561 2 554 1 INV1S $T=324880 467160 1 180 $X=323640 $Y=466780
X536 562 2 530 1 INV1S $T=324880 497400 1 180 $X=323640 $Y=497020
X537 540 2 553 1 INV1S $T=324880 517560 1 180 $X=323640 $Y=517180
X538 566 2 540 1 INV1S $T=326120 517560 1 180 $X=324880 $Y=517180
X539 579 2 580 1 INV1S $T=329220 467160 0 0 $X=329220 $Y=466780
X540 574 2 586 1 INV1S $T=334180 467160 0 180 $X=332940 $Y=461740
X541 560 2 573 1 INV1S $T=334800 457080 1 180 $X=333560 $Y=456700
X542 565 2 588 1 INV1S $T=334800 467160 1 180 $X=333560 $Y=466780
X543 600 2 595 1 INV1S $T=336660 497400 0 180 $X=335420 $Y=491980
X544 606 2 575 1 INV1S $T=337280 517560 1 180 $X=336040 $Y=517180
X545 589 2 603 1 INV1S $T=338520 487320 1 180 $X=337280 $Y=486940
X546 632 2 629 1 INV1S $T=344100 477240 1 180 $X=342860 $Y=476860
X547 642 2 621 1 INV1S $T=345960 477240 1 180 $X=344720 $Y=476860
X548 612 2 628 1 INV1S $T=344720 517560 0 0 $X=344720 $Y=517180
X549 35 2 654 1 INV1S $T=347820 537720 0 0 $X=347820 $Y=537340
X550 659 2 653 1 INV1S $T=349680 447000 1 180 $X=348440 $Y=446620
X551 607 2 648 1 INV1S $T=349680 507480 0 180 $X=348440 $Y=502060
X552 593 2 662 1 INV1S $T=349060 537720 0 0 $X=349060 $Y=537340
X553 668 2 656 1 INV1S $T=351540 436920 0 0 $X=351540 $Y=436540
X554 674 2 667 1 INV1S $T=352780 487320 1 180 $X=351540 $Y=486940
X555 660 2 661 1 INV1S $T=352780 497400 1 180 $X=351540 $Y=497020
X556 657 2 658 1 INV1S $T=354640 497400 0 180 $X=353400 $Y=491980
X557 647 2 672 1 INV1S $T=355880 517560 1 180 $X=354640 $Y=517180
X558 707 2 705 1 INV1S $T=362080 467160 0 180 $X=360840 $Y=461740
X559 37 2 709 1 INV1S $T=360840 537720 0 0 $X=360840 $Y=537340
X560 715 2 711 1 INV1S $T=363940 447000 1 180 $X=362700 $Y=446620
X561 732 2 710 1 INV1S $T=365180 447000 1 180 $X=363940 $Y=446620
X562 688 2 721 1 INV1S $T=365180 426840 0 0 $X=365180 $Y=426460
X563 727 2 719 1 INV1S $T=366420 517560 0 180 $X=365180 $Y=512140
X564 742 2 718 1 INV1S $T=368900 426840 1 180 $X=367660 $Y=426460
X565 40 2 746 1 INV1S $T=368280 537720 0 0 $X=368280 $Y=537340
X566 736 2 741 1 INV1S $T=370140 467160 1 180 $X=368900 $Y=466780
X567 722 2 747 1 INV1S $T=370760 487320 0 180 $X=369520 $Y=481900
X568 41 2 752 1 INV1S $T=369520 537720 0 0 $X=369520 $Y=537340
X569 761 2 757 1 INV1S $T=372620 477240 1 180 $X=371380 $Y=476860
X570 759 2 760 1 INV1S $T=372000 457080 1 0 $X=372000 $Y=451660
X571 731 2 749 1 INV1S $T=375100 436920 0 180 $X=373860 $Y=431500
X572 782 2 778 1 INV1S $T=378200 467160 1 180 $X=376960 $Y=466780
X573 755 2 769 1 INV1S $T=377580 517560 0 0 $X=377580 $Y=517180
X574 802 2 762 1 INV1S $T=380060 467160 1 180 $X=378820 $Y=466780
X575 803 2 797 1 INV1S $T=381920 457080 0 180 $X=380680 $Y=451660
X576 776 2 792 1 INV1S $T=383160 497400 0 180 $X=381920 $Y=491980
X577 42 2 813 1 INV1S $T=381920 537720 0 0 $X=381920 $Y=537340
X578 806 2 767 1 INV1S $T=382540 477240 1 0 $X=382540 $Y=471820
X579 43 2 820 1 INV1S $T=383160 537720 0 0 $X=383160 $Y=537340
X580 822 2 819 1 INV1S $T=385020 477240 0 180 $X=383780 $Y=471820
X581 795 2 777 1 INV1S $T=385020 497400 0 180 $X=383780 $Y=491980
X582 781 2 798 1 INV1S $T=385020 507480 1 180 $X=383780 $Y=507100
X583 826 2 796 1 INV1S $T=385640 436920 1 180 $X=384400 $Y=436540
X584 815 2 823 1 INV1S $T=385640 477240 1 180 $X=384400 $Y=476860
X585 832 2 837 1 INV1S $T=388740 457080 1 180 $X=387500 $Y=456700
X586 802 2 827 1 INV1S $T=387500 467160 0 0 $X=387500 $Y=466780
X587 825 2 835 1 INV1S $T=388740 487320 1 180 $X=387500 $Y=486940
X588 847 2 841 1 INV1S $T=388740 497400 1 180 $X=387500 $Y=497020
X589 754 2 785 1 INV1S $T=388740 527640 0 180 $X=387500 $Y=522220
X590 828 2 854 1 INV1S $T=389360 457080 1 0 $X=389360 $Y=451660
X591 877 2 829 1 INV1S $T=391220 457080 1 180 $X=389980 $Y=456700
X592 867 2 856 1 INV1S $T=393080 517560 1 180 $X=391840 $Y=517180
X593 864 2 802 1 INV1S $T=393700 467160 1 180 $X=392460 $Y=466780
X594 866 2 860 1 INV1S $T=394940 507480 1 180 $X=393700 $Y=507100
X595 858 2 852 1 INV1S $T=395560 497400 0 180 $X=394320 $Y=491980
X596 858 2 839 1 INV1S $T=395560 507480 0 180 $X=394320 $Y=502060
X597 874 2 863 1 INV1S $T=396180 457080 0 180 $X=394940 $Y=451660
X598 858 2 870 1 INV1S $T=394940 467160 0 0 $X=394940 $Y=466780
X599 869 2 868 1 INV1S $T=397420 436920 1 180 $X=396180 $Y=436540
X600 891 2 861 1 INV1S $T=398660 436920 1 180 $X=397420 $Y=436540
X601 882 2 857 1 INV1S $T=398660 497400 1 180 $X=397420 $Y=497020
X602 806 2 766 1 INV1S $T=401760 457080 1 180 $X=400520 $Y=456700
X603 929 2 905 1 INV1S $T=406100 507480 0 180 $X=404860 $Y=502060
X604 931 2 52 1 INV1S $T=407340 406680 0 0 $X=407340 $Y=406300
X605 940 2 938 1 INV1S $T=409820 426840 1 180 $X=408580 $Y=426460
X606 948 2 951 1 INV1S $T=411680 467160 0 180 $X=410440 $Y=461740
X607 942 2 957 1 INV1S $T=411060 487320 0 0 $X=411060 $Y=486940
X608 946 2 906 1 INV1S $T=412300 527640 1 0 $X=412300 $Y=522220
X609 936 2 937 1 INV1S $T=412920 447000 1 0 $X=412920 $Y=441580
X610 988 2 54 1 INV1S $T=420980 426840 0 180 $X=419740 $Y=421420
X611 984 2 894 1 INV1S $T=422220 447000 0 0 $X=422220 $Y=446620
X612 1001 2 999 1 INV1S $T=427180 447000 0 180 $X=425940 $Y=441580
X613 1006 2 917 1 INV1S $T=427180 477240 1 180 $X=425940 $Y=476860
X614 858 2 1017 1 INV1S $T=427800 467160 0 0 $X=427800 $Y=466780
X615 1015 2 994 1 INV1S $T=429040 537720 1 180 $X=427800 $Y=537340
X616 1009 2 1012 1 INV1S $T=429660 477240 1 180 $X=428420 $Y=476860
X617 1022 2 1016 1 INV1S $T=430280 436920 0 180 $X=429040 $Y=431500
X618 59 2 62 1 INV1S $T=430280 537720 0 0 $X=430280 $Y=537340
X619 1014 2 1027 1 INV1S $T=432760 497400 0 0 $X=432760 $Y=497020
X620 1049 2 1006 1 INV1S $T=436480 497400 0 180 $X=435240 $Y=491980
X621 1047 2 753 1 INV1S $T=437100 457080 1 180 $X=435860 $Y=456700
X622 916 2 1025 1 INV1S $T=437100 507480 1 180 $X=435860 $Y=507100
X623 1004 2 1053 1 INV1S $T=437100 487320 1 0 $X=437100 $Y=481900
X624 1034 2 63 1 INV1S $T=437100 527640 0 0 $X=437100 $Y=527260
X625 1006 2 1059 1 INV1S $T=437720 497400 1 0 $X=437720 $Y=491980
X626 993 2 1038 1 INV1S $T=440200 467160 0 180 $X=438960 $Y=461740
X627 1063 2 1052 1 INV1S $T=440820 436920 1 180 $X=439580 $Y=436540
X628 1031 2 1056 1 INV1S $T=441440 436920 0 180 $X=440200 $Y=431500
X629 1039 2 1070 1 INV1S $T=443300 467160 1 180 $X=442060 $Y=466780
X630 65 2 989 1 INV1S $T=442680 497400 0 0 $X=442680 $Y=497020
X631 858 2 1079 1 INV1S $T=443920 467160 0 0 $X=443920 $Y=466780
X632 1087 2 1058 1 INV1S $T=445160 537720 1 180 $X=443920 $Y=537340
X633 1080 2 1076 1 INV1S $T=445160 416760 1 0 $X=445160 $Y=411340
X634 1037 2 67 1 INV1S $T=445160 426840 0 0 $X=445160 $Y=426460
X635 1039 2 1095 1 INV1S $T=445780 467160 0 0 $X=445780 $Y=466780
X636 1069 2 1096 1 INV1S $T=445780 487320 0 0 $X=445780 $Y=486940
X637 1047 2 1104 1 INV1S $T=446400 457080 0 0 $X=446400 $Y=456700
X638 1093 2 1107 1 INV1S $T=449500 507480 1 0 $X=449500 $Y=502060
X639 1101 2 1118 1 INV1S $T=451360 477240 1 0 $X=451360 $Y=471820
X640 1135 2 1120 1 INV1S $T=454460 406680 1 180 $X=453220 $Y=406300
X641 1024 2 1023 1 INV1S $T=454460 497400 1 180 $X=453220 $Y=497020
X642 1123 2 1119 1 INV1S $T=455080 517560 0 180 $X=453840 $Y=512140
X643 1092 2 72 1 INV1S $T=455700 436920 0 180 $X=454460 $Y=431500
X644 1130 2 1134 1 INV1S $T=454460 507480 0 0 $X=454460 $Y=507100
X645 1108 2 1139 1 INV1S $T=455700 467160 1 0 $X=455700 $Y=461740
X646 1059 2 1121 1 INV1S $T=456940 497400 1 180 $X=455700 $Y=497020
X647 1126 2 1128 1 INV1S $T=457560 457080 0 180 $X=456320 $Y=451660
X648 1110 2 1151 1 INV1S $T=458180 497400 0 0 $X=458180 $Y=497020
X649 1159 2 69 1 INV1S $T=460040 537720 1 180 $X=458800 $Y=537340
X650 1143 2 1160 1 INV1S $T=460660 406680 1 0 $X=460660 $Y=401260
X651 1170 2 53 1 INV1S $T=463760 487320 1 180 $X=462520 $Y=486940
X652 1157 2 1176 1 INV1S $T=463140 497400 0 0 $X=463140 $Y=497020
X653 1174 2 1180 1 INV1S $T=463760 487320 0 0 $X=463760 $Y=486940
X654 1167 2 1177 1 INV1S $T=463760 507480 1 0 $X=463760 $Y=502060
X655 1141 2 1187 1 INV1S $T=465620 467160 0 0 $X=465620 $Y=466780
X656 1192 2 1203 1 INV1S $T=468720 406680 1 0 $X=468720 $Y=401260
X657 1196 2 1169 1 INV1S $T=468720 416760 1 0 $X=468720 $Y=411340
X658 1189 2 1204 1 INV1S $T=468720 447000 1 0 $X=468720 $Y=441580
X659 1195 2 1201 1 INV1S $T=468720 497400 1 0 $X=468720 $Y=491980
X660 1211 2 1173 1 INV1S $T=472440 416760 1 180 $X=471200 $Y=416380
X661 1229 2 1216 1 INV1S $T=476160 507480 0 180 $X=474920 $Y=502060
X662 1182 2 1225 1 INV1S $T=476160 477240 1 0 $X=476160 $Y=471820
X663 1193 2 1226 1 INV1S $T=479880 447000 1 180 $X=478640 $Y=446620
X664 1224 2 1242 1 INV1S $T=479880 457080 0 0 $X=479880 $Y=456700
X665 1251 2 1222 1 INV1S $T=481740 416760 0 180 $X=480500 $Y=411340
X666 1234 2 1256 1 INV1S $T=481740 467160 1 0 $X=481740 $Y=461740
X667 92 2 86 1 INV1S $T=482980 537720 1 180 $X=481740 $Y=537340
X668 1244 2 1263 1 INV1S $T=485460 467160 0 0 $X=485460 $Y=466780
X669 1258 2 1230 1 INV1S $T=486080 426840 1 0 $X=486080 $Y=421420
X670 1235 2 1255 1 INV1S $T=486080 487320 0 0 $X=486080 $Y=486940
X671 1245 2 1264 1 INV1S $T=487320 467160 1 0 $X=487320 $Y=461740
X672 1265 2 1268 1 INV1S $T=487940 447000 1 0 $X=487940 $Y=441580
X673 1273 2 1257 1 INV1S $T=491040 426840 0 180 $X=489800 $Y=421420
X674 1290 2 1261 1 INV1S $T=497240 416760 0 180 $X=496000 $Y=411340
X675 1292 2 1284 1 INV1S $T=499100 416760 1 180 $X=497860 $Y=416380
X676 1299 2 1285 1 INV1S $T=500960 457080 0 180 $X=499720 $Y=451660
X677 1302 2 1283 1 INV1S $T=503440 457080 0 180 $X=502200 $Y=451660
X678 1276 2 1300 1 INV1S $T=502200 467160 0 0 $X=502200 $Y=466780
X679 1304 2 1301 1 INV1S $T=504060 447000 1 0 $X=504060 $Y=441580
X680 1303 2 1296 1 INV1S $T=504680 487320 1 0 $X=504680 $Y=481900
X681 1321 2 1295 1 INV1S $T=508400 436920 0 180 $X=507160 $Y=431500
X682 104 2 94 1 INV1S $T=507160 537720 0 0 $X=507160 $Y=537340
X683 1316 2 102 1 INV1S $T=508400 527640 1 0 $X=508400 $Y=522220
X684 1319 2 99 1 INV1S $T=511500 527640 1 180 $X=510260 $Y=527260
X685 1325 2 1272 1 INV1S $T=510880 416760 1 0 $X=510880 $Y=411340
X686 1350 2 1320 1 INV1S $T=513360 436920 1 180 $X=512120 $Y=436540
X687 1351 2 1314 1 INV1S $T=516460 467160 0 180 $X=515220 $Y=461740
X688 1343 2 111 1 INV1S $T=517700 477240 0 180 $X=516460 $Y=471820
X689 1344 2 1334 1 INV1S $T=519560 497400 0 180 $X=518320 $Y=491980
X690 1338 2 100 1 INV1S $T=518940 507480 0 0 $X=518940 $Y=507100
X691 1348 2 110 1 INV1S $T=520800 457080 0 180 $X=519560 $Y=451660
X692 1339 2 1327 1 INV1S $T=519560 487320 1 0 $X=519560 $Y=481900
X693 117 2 1305 1 INV1S $T=520800 517560 0 180 $X=519560 $Y=512140
X694 1347 2 107 1 INV1S $T=521420 527640 0 180 $X=520180 $Y=522220
X695 1349 2 1330 1 INV1S $T=522040 416760 1 180 $X=520800 $Y=416380
X696 1341 2 1315 1 INV1S $T=522040 507480 1 0 $X=522040 $Y=502060
X697 1358 2 1355 1 INV1S $T=524520 406680 0 180 $X=523280 $Y=401260
X698 1379 2 1346 1 INV1S $T=530720 436920 0 180 $X=529480 $Y=431500
X699 1388 2 1372 1 INV1S $T=533200 457080 0 180 $X=531960 $Y=451660
X700 1380 2 129 1 INV1S $T=533820 537720 1 180 $X=532580 $Y=537340
X701 1392 2 118 1 INV1S $T=533820 527640 0 0 $X=533820 $Y=527260
X702 1396 2 1394 1 INV1S $T=535680 396600 1 180 $X=534440 $Y=396220
X703 135 2 139 1 INV1S $T=540020 396600 1 0 $X=540020 $Y=391180
X704 1385 2 1425 1 INV1S $T=543120 477240 1 180 $X=541880 $Y=476860
X705 1426 2 126 1 INV1S $T=541880 537720 0 0 $X=541880 $Y=537340
X706 1395 2 1432 1 INV1S $T=543120 406680 1 0 $X=543120 $Y=401260
X707 1399 2 1441 1 INV1S $T=543740 457080 0 0 $X=543740 $Y=456700
X708 1431 2 119 1 INV1S $T=544980 527640 1 180 $X=543740 $Y=527260
X709 1429 2 1435 1 INV1S $T=544360 396600 1 0 $X=544360 $Y=391180
X710 1421 2 1440 1 INV1S $T=545600 406680 1 0 $X=545600 $Y=401260
X711 1442 2 1449 1 INV1S $T=547460 416760 1 0 $X=547460 $Y=411340
X712 1444 2 1433 1 INV1S $T=550560 477240 0 0 $X=550560 $Y=476860
X713 1437 2 1454 1 INV1S $T=553040 487320 1 180 $X=551800 $Y=486940
X714 1455 2 1459 1 INV1S $T=553660 406680 1 180 $X=552420 $Y=406300
X715 117 2 154 1 INV1S $T=555520 537720 0 0 $X=555520 $Y=537340
X716 1478 2 1484 1 INV1S $T=557380 406680 1 0 $X=557380 $Y=401260
X717 1489 2 1476 1 INV1S $T=558620 436920 1 180 $X=557380 $Y=436540
X718 1482 2 1470 1 INV1S $T=558620 447000 1 180 $X=557380 $Y=446620
X719 1438 2 1472 1 INV1S $T=558000 507480 1 0 $X=558000 $Y=502060
X720 1450 2 1492 1 INV1S $T=558620 457080 0 0 $X=558620 $Y=456700
X721 1494 2 1501 1 INV1S $T=561720 487320 0 0 $X=561720 $Y=486940
X722 1485 2 1515 1 INV1S $T=563580 416760 1 0 $X=563580 $Y=411340
X723 1502 2 1511 1 INV1S $T=565440 406680 1 0 $X=565440 $Y=401260
X724 1505 2 1527 1 INV1S $T=566680 426840 1 0 $X=566680 $Y=421420
X725 1529 2 1520 1 INV1S $T=569160 436920 1 0 $X=569160 $Y=431500
X726 1526 2 1539 1 INV1S $T=569780 457080 0 0 $X=569780 $Y=456700
X727 1533 2 1552 1 INV1S $T=572880 447000 0 0 $X=572880 $Y=446620
X728 1545 2 1294 1 INV1S $T=572880 537720 1 0 $X=572880 $Y=532300
X729 1413 2 1538 1 INV1S $T=573500 487320 1 0 $X=573500 $Y=481900
X730 1560 2 1537 1 INV1S $T=575360 507480 0 180 $X=574120 $Y=502060
X731 1427 2 1569 1 INV1S $T=575360 396600 1 0 $X=575360 $Y=391180
X732 1547 2 1564 1 INV1S $T=575360 426840 1 0 $X=575360 $Y=421420
X733 1573 2 1562 1 INV1S $T=577840 507480 0 180 $X=576600 $Y=502060
X734 1554 2 1567 1 INV1S $T=578460 416760 0 180 $X=577220 $Y=411340
X735 1593 2 1615 1 INV1S $T=582180 396600 0 0 $X=582180 $Y=396220
X736 1503 2 1585 1 INV1S $T=585900 406680 1 180 $X=584660 $Y=406300
X737 1503 2 1613 1 INV1S $T=585900 416760 0 0 $X=585900 $Y=416380
X738 1581 2 1622 1 INV1S $T=586520 487320 1 0 $X=586520 $Y=481900
X739 1607 2 1360 1 INV1S $T=586520 537720 1 0 $X=586520 $Y=532300
X740 1599 2 1627 1 INV1S $T=587140 527640 1 0 $X=587140 $Y=522220
X741 1589 2 1603 1 INV1S $T=589000 406680 1 0 $X=589000 $Y=401260
X742 1572 2 1605 1 INV1S $T=589000 447000 1 0 $X=589000 $Y=441580
X743 1568 2 1641 1 INV1S $T=590860 517560 1 0 $X=590860 $Y=512140
X744 1597 2 1618 1 INV1S $T=591480 406680 0 0 $X=591480 $Y=406300
X745 1616 2 1625 1 INV1S $T=592720 416760 1 180 $X=591480 $Y=416380
X746 1523 2 1633 1 INV1S $T=592100 507480 1 0 $X=592100 $Y=502060
X747 1621 2 1637 1 INV1S $T=594580 477240 1 0 $X=594580 $Y=471820
X748 1600 2 1651 1 INV1S $T=594580 527640 1 0 $X=594580 $Y=522220
X749 1361 2 1660 1 INV1S $T=598300 406680 0 0 $X=598300 $Y=406300
X750 1612 2 1668 1 INV1S $T=599540 517560 1 0 $X=599540 $Y=512140
X751 1664 2 1667 1 INV1S $T=599540 527640 1 0 $X=599540 $Y=522220
X752 1566 2 1701 1 INV1S $T=601400 477240 0 0 $X=601400 $Y=476860
X753 1661 2 1694 1 INV1S $T=602640 467160 1 0 $X=602640 $Y=461740
X754 1588 2 1692 1 INV1S $T=603880 467160 0 0 $X=603880 $Y=466780
X755 1517 2 1691 1 INV1S $T=605120 487320 1 0 $X=605120 $Y=481900
X756 1671 2 1679 1 INV1S $T=606980 527640 1 180 $X=605740 $Y=527260
X757 1659 2 1704 1 INV1S $T=606980 507480 1 0 $X=606980 $Y=502060
X758 1570 2 1716 1 INV1S $T=608220 416760 0 0 $X=608220 $Y=416380
X759 1657 2 1703 1 INV1S $T=608220 527640 1 0 $X=608220 $Y=522220
X760 1630 2 1719 1 INV1S $T=611940 507480 0 0 $X=611940 $Y=507100
X761 1592 2 1733 1 INV1S $T=616280 447000 0 0 $X=616280 $Y=446620
X762 1662 2 1741 1 INV1S $T=617520 416760 1 0 $X=617520 $Y=411340
X763 1528 2 1728 1 INV1S $T=618760 447000 0 0 $X=618760 $Y=446620
X764 1722 2 1744 1 INV1S $T=619380 527640 1 0 $X=619380 $Y=522220
X765 1683 2 1749 1 INV1S $T=620000 517560 1 0 $X=620000 $Y=512140
X766 1700 2 1750 1 INV1S $T=621860 436920 0 0 $X=621860 $Y=436540
X767 1740 2 188 1 INV1S $T=623100 537720 1 0 $X=623100 $Y=532300
X768 1565 2 1748 1 INV1S $T=623720 477240 1 0 $X=623720 $Y=471820
X769 1662 2 1763 1 INV1S $T=625580 416760 1 0 $X=625580 $Y=411340
X770 1718 2 1792 1 INV1S $T=626820 447000 0 0 $X=626820 $Y=446620
X771 1735 2 1769 1 INV1S $T=628060 416760 0 0 $X=628060 $Y=416380
X772 1678 2 1781 1 INV1S $T=629300 426840 1 0 $X=629300 $Y=421420
X773 1772 2 1777 1 INV1S $T=629920 487320 1 0 $X=629920 $Y=481900
X774 1757 2 1778 1 INV1S $T=631160 436920 1 0 $X=631160 $Y=431500
X775 1756 2 1782 1 INV1S $T=632400 517560 0 180 $X=631160 $Y=512140
X776 1761 2 1794 1 INV1S $T=633020 497400 1 0 $X=633020 $Y=491980
X777 1775 2 1799 1 INV1S $T=635500 487320 1 0 $X=635500 $Y=481900
X778 193 2 1801 1 INV1S $T=637360 396600 0 0 $X=637360 $Y=396220
X779 1422 2 197 1 INV1S $T=639220 527640 1 0 $X=639220 $Y=522220
X780 1784 2 1821 1 INV1S $T=641700 487320 0 0 $X=641700 $Y=486940
X781 191 2 1825 1 INV1S $T=642320 396600 1 0 $X=642320 $Y=391180
X782 1745 2 199 1 INV1S $T=642940 537720 1 0 $X=642940 $Y=532300
X783 1830 2 1832 1 INV1S $T=643560 436920 0 0 $X=643560 $Y=436540
X784 1407 2 200 1 INV1S $T=645420 517560 1 0 $X=645420 $Y=512140
X785 1617 2 201 1 INV1S $T=645420 527640 0 0 $X=645420 $Y=527260
X786 1822 2 1845 1 INV1S $T=646040 396600 1 0 $X=646040 $Y=391180
X787 1826 2 1847 1 INV1S $T=646040 467160 1 0 $X=646040 $Y=461740
X788 1843 2 178 1 INV1S $T=647900 537720 0 0 $X=647900 $Y=537340
X789 1834 2 1854 1 INV1S $T=648520 416760 0 0 $X=648520 $Y=416380
X790 1841 2 1851 1 INV1S $T=649760 467160 0 180 $X=648520 $Y=461740
X791 1809 2 1873 1 INV1S $T=652240 457080 1 0 $X=652240 $Y=451660
X792 1881 2 1856 1 INV1S $T=656580 537720 0 180 $X=655340 $Y=532300
X793 1883 2 1840 1 INV1S $T=660920 517560 0 180 $X=659680 $Y=512140
X794 1687 2 221 1 INV1S $T=660300 537720 1 0 $X=660300 $Y=532300
X795 1903 2 1861 1 INV1S $T=662160 527640 1 180 $X=660920 $Y=527260
X796 1887 2 1860 1 INV1S $T=664020 517560 0 180 $X=662780 $Y=512140
X797 1889 2 1902 1 INV1S $T=667120 426840 1 0 $X=667120 $Y=421420
X798 1915 2 1911 1 INV1S $T=672080 416760 1 180 $X=670840 $Y=416380
X799 1780 2 1941 1 INV1S $T=670840 527640 1 0 $X=670840 $Y=522220
X800 1899 2 1923 1 INV1S $T=675180 436920 0 180 $X=673940 $Y=431500
X801 1932 2 1926 1 INV1S $T=676420 457080 1 180 $X=675180 $Y=456700
X802 1928 2 1933 1 INV1S $T=675800 447000 1 0 $X=675800 $Y=441580
X803 1908 2 1931 1 INV1S $T=675800 447000 0 0 $X=675800 $Y=446620
X804 1918 2 1944 1 INV1S $T=677660 416760 1 0 $X=677660 $Y=411340
X805 1951 2 1943 1 INV1S $T=680140 487320 0 180 $X=678900 $Y=481900
X806 1935 2 1920 1 INV1S $T=681380 537720 0 180 $X=680140 $Y=532300
X807 1953 2 1948 1 INV1S $T=680760 426840 0 0 $X=680760 $Y=426460
X808 1902 2 1959 1 INV1S $T=682000 426840 1 0 $X=682000 $Y=421420
X809 1957 2 1965 1 INV1S $T=682000 467160 0 0 $X=682000 $Y=466780
X810 1904 2 249 1 INV1S $T=682620 396600 0 0 $X=682620 $Y=396220
X811 1961 2 1970 1 INV1S $T=685100 436920 0 0 $X=685100 $Y=436540
X812 1955 2 1989 1 INV1S $T=688820 406680 1 0 $X=688820 $Y=401260
X813 1931 2 1966 1 INV1S $T=690680 447000 1 180 $X=689440 $Y=446620
X814 1939 2 1991 1 INV1S $T=690060 436920 1 0 $X=690060 $Y=431500
X815 1931 2 1994 1 INV1S $T=690680 447000 0 0 $X=690680 $Y=446620
X816 258 2 1982 1 INV1S $T=690680 537720 0 0 $X=690680 $Y=537340
X817 1998 2 2005 1 INV1S $T=692540 487320 0 0 $X=692540 $Y=486940
X818 2000 2 2006 1 INV1S $T=692540 497400 0 0 $X=692540 $Y=497020
X819 1988 2 2023 1 INV1S $T=694400 477240 1 0 $X=694400 $Y=471820
X820 256 2 2034 1 INV1S $T=696260 447000 1 0 $X=696260 $Y=441580
X821 1978 2 2025 1 INV1S $T=696880 457080 1 0 $X=696880 $Y=451660
X822 2028 2 2041 1 INV1S $T=698120 457080 1 0 $X=698120 $Y=451660
X823 2054 2 2018 1 INV1S $T=699980 487320 1 180 $X=698740 $Y=486940
X824 2027 2 2035 1 INV1S $T=702460 497400 1 180 $X=701220 $Y=497020
X825 1916 2 2057 1 INV1S $T=705560 477240 1 180 $X=704320 $Y=476860
X826 1946 2 2073 1 INV1S $T=704320 527640 1 0 $X=704320 $Y=522220
X827 2048 2 2087 1 INV1S $T=706800 497400 1 0 $X=706800 $Y=491980
X828 2069 2 2089 1 INV1S $T=707420 406680 1 0 $X=707420 $Y=401260
X829 2076 2 2091 1 INV1S $T=707420 426840 1 0 $X=707420 $Y=421420
X830 2077 2 2079 1 INV1S $T=709280 416760 1 180 $X=708040 $Y=416380
X831 2075 2 2084 1 INV1S $T=709900 396600 1 180 $X=708660 $Y=396220
X832 2103 2 2096 1 INV1S $T=711760 497400 0 180 $X=710520 $Y=491980
X833 2111 2 2114 1 INV1S $T=712380 416760 1 0 $X=712380 $Y=411340
X834 2092 2 2119 1 INV1S $T=712380 477240 0 0 $X=712380 $Y=476860
X835 2114 2 2133 1 INV1S $T=714240 406680 1 0 $X=714240 $Y=401260
X836 2011 2 2140 1 INV1S $T=715480 487320 0 0 $X=715480 $Y=486940
X837 2063 2 2137 1 INV1S $T=717960 447000 0 180 $X=716720 $Y=441580
X838 2126 2 2141 1 INV1S $T=717960 497400 0 180 $X=716720 $Y=491980
X839 2107 2 2104 1 INV1S $T=717340 477240 0 0 $X=717340 $Y=476860
X840 278 2 2108 1 INV1S $T=718580 537720 1 180 $X=717340 $Y=537340
X841 2129 2 2163 1 INV1S $T=717960 436920 1 0 $X=717960 $Y=431500
X842 2123 2 2157 1 INV1S $T=719200 527640 0 0 $X=719200 $Y=527260
X843 2152 2 2160 1 INV1S $T=719820 426840 1 0 $X=719820 $Y=421420
X844 2068 2 2155 1 INV1S $T=719820 467160 0 0 $X=719820 $Y=466780
X845 2121 2 2166 1 INV1S $T=720440 416760 1 0 $X=720440 $Y=411340
X846 279 2 2162 1 INV1S $T=720440 537720 0 0 $X=720440 $Y=537340
X847 2158 2 2171 1 INV1S $T=722920 487320 0 0 $X=722920 $Y=486940
X848 2153 2 2161 1 INV1S $T=724780 457080 0 180 $X=723540 $Y=451660
X849 280 2 2173 1 INV1S $T=724160 396600 0 0 $X=724160 $Y=396220
X850 2146 2 2168 1 INV1S $T=725400 406680 1 180 $X=724160 $Y=406300
X851 2132 2 2182 1 INV1S $T=724160 487320 0 0 $X=724160 $Y=486940
X852 2167 2 2187 1 INV1S $T=724780 497400 1 0 $X=724780 $Y=491980
X853 283 2 2178 1 INV1S $T=726640 537720 1 180 $X=725400 $Y=537340
X854 2184 2 2193 1 INV1S $T=726640 457080 0 0 $X=726640 $Y=456700
X855 2177 2 2212 1 INV1S $T=728500 527640 0 0 $X=728500 $Y=527260
X856 2001 2 2214 1 INV1S $T=729120 396600 1 0 $X=729120 $Y=391180
X857 1976 2 2206 1 INV1S $T=730360 457080 1 0 $X=730360 $Y=451660
X858 2021 2 2223 1 INV1S $T=730980 467160 1 0 $X=730980 $Y=461740
X859 2060 2 2222 1 INV1S $T=732220 457080 0 0 $X=732220 $Y=456700
X860 2217 2 2227 1 INV1S $T=732840 527640 1 0 $X=732840 $Y=522220
X861 2039 2 2238 1 INV1S $T=735320 416760 1 0 $X=735320 $Y=411340
X862 2242 2 2246 1 INV1S $T=736560 416760 1 0 $X=736560 $Y=411340
X863 2241 2 2247 1 INV1S $T=738420 497400 0 180 $X=737180 $Y=491980
X864 2226 2 2265 1 INV1S $T=740900 477240 0 0 $X=740900 $Y=476860
X865 2253 2 2266 1 INV1S $T=740900 527640 0 0 $X=740900 $Y=527260
X866 2210 2 2277 1 INV1S $T=741520 426840 0 0 $X=741520 $Y=426460
X867 2236 2 2287 1 INV1S $T=744000 487320 0 0 $X=744000 $Y=486940
X868 2245 2 2308 1 INV1S $T=750200 457080 0 180 $X=748960 $Y=451660
X869 2254 2 2313 1 INV1S $T=749580 457080 0 0 $X=749580 $Y=456700
X870 2250 2 2310 1 INV1S $T=750820 517560 1 180 $X=749580 $Y=517180
X871 1995 2 2292 1 INV1S $T=750200 406680 0 0 $X=750200 $Y=406300
X872 2245 2 2336 1 INV1S $T=750820 457080 0 0 $X=750820 $Y=456700
X873 2325 2 2322 1 INV1S $T=753300 477240 1 180 $X=752060 $Y=476860
X874 294 2 293 1 INV1S $T=753920 537720 1 180 $X=752680 $Y=537340
X875 2264 2 2331 1 INV1S $T=753300 467160 0 0 $X=753300 $Y=466780
X876 2273 2 2335 1 INV1S $T=753920 527640 1 0 $X=753920 $Y=522220
X877 2260 2 2361 1 INV1S $T=761360 426840 1 180 $X=760120 $Y=426460
X878 2280 2 2348 1 INV1S $T=760120 527640 1 0 $X=760120 $Y=522220
X879 2272 2 2370 1 INV1S $T=761980 426840 1 0 $X=761980 $Y=421420
X880 2357 2 2377 1 INV1S $T=765080 517560 0 180 $X=763840 $Y=512140
X881 2244 2 2362 1 INV1S $T=764460 436920 0 0 $X=764460 $Y=436540
X882 2305 2 2392 1 INV1S $T=765700 517560 0 0 $X=765700 $Y=517180
X883 2390 2 2389 1 INV1S $T=766320 537720 1 0 $X=766320 $Y=532300
X884 2368 2 2395 1 INV1S $T=766940 457080 0 0 $X=766940 $Y=456700
X885 2318 2 2406 1 INV1S $T=767560 517560 0 0 $X=767560 $Y=517180
X886 2375 2 2413 1 INV1S $T=768180 527640 0 0 $X=768180 $Y=527260
X887 2399 2 2411 1 INV1S $T=768800 507480 1 0 $X=768800 $Y=502060
X888 2402 2 2414 1 INV1S $T=770660 457080 1 0 $X=770660 $Y=451660
X889 2403 2 2409 1 INV1S $T=770660 537720 0 0 $X=770660 $Y=537340
X890 298 2 2419 1 INV1S $T=772520 396600 1 0 $X=772520 $Y=391180
X891 2383 2 2431 1 INV1S $T=773760 447000 0 0 $X=773760 $Y=446620
X892 303 2 2424 1 INV1S $T=774380 396600 0 0 $X=774380 $Y=396220
X893 302 2 2439 1 INV1S $T=776860 396600 0 0 $X=776860 $Y=396220
X894 2428 2 2444 1 INV1S $T=777480 487320 0 0 $X=777480 $Y=486940
X895 2365 2 2412 1 INV1S $T=777480 517560 1 0 $X=777480 $Y=512140
X896 2364 2 2441 1 INV1S $T=779960 517560 0 180 $X=778720 $Y=512140
X897 2391 2 2454 1 INV1S $T=779960 517560 1 0 $X=779960 $Y=512140
X898 2450 2 2456 1 INV1S $T=783060 436920 0 180 $X=781820 $Y=431500
X899 309 2 2471 1 INV1S $T=783680 537720 0 0 $X=783680 $Y=537340
X900 2458 2 2481 1 INV1S $T=784300 426840 0 0 $X=784300 $Y=426460
X901 2387 2 2482 1 INV1S $T=785540 507480 0 0 $X=785540 $Y=507100
X902 315 2 2496 1 INV1S $T=792360 537720 0 0 $X=792360 $Y=537340
X903 2512 2 2524 1 INV1S $T=799180 477240 0 0 $X=799180 $Y=476860
X904 2522 2 2534 1 INV1S $T=801040 477240 0 0 $X=801040 $Y=476860
X905 2530 2 2562 1 INV1S $T=807860 477240 1 0 $X=807860 $Y=471820
X906 2539 2 2556 1 INV1S $T=811580 487320 0 180 $X=810340 $Y=481900
X907 2575 2 2599 1 INV1S $T=814680 447000 1 0 $X=814680 $Y=441580
X908 2582 2 2584 1 INV1S $T=815920 467160 0 180 $X=814680 $Y=461740
X909 2542 2 2591 1 INV1S $T=815920 487320 1 0 $X=815920 $Y=481900
X910 2505 2 2592 1 INV1S $T=815920 487320 0 0 $X=815920 $Y=486940
X911 2595 2 2589 1 INV1S $T=818400 426840 0 180 $X=817160 $Y=421420
X912 2570 2 2597 1 INV1S $T=817160 467160 0 0 $X=817160 $Y=466780
X913 2568 2 2609 1 INV1S $T=818400 487320 1 0 $X=818400 $Y=481900
X914 2561 2 2605 1 INV1S $T=819640 467160 1 0 $X=819640 $Y=461740
X915 2612 2 2616 1 INV1S $T=820880 467160 0 0 $X=820880 $Y=466780
X916 2564 2 2633 1 INV1S $T=822120 426840 0 0 $X=822120 $Y=426460
X917 2571 2 2620 1 INV1S $T=822740 467160 1 0 $X=822740 $Y=461740
X918 2625 2 2630 1 INV1S $T=823980 416760 0 0 $X=823980 $Y=416380
X919 2567 2 2636 1 INV1S $T=824600 436920 0 0 $X=824600 $Y=436540
X920 2600 2 2637 1 INV1S $T=825220 457080 1 0 $X=825220 $Y=451660
X921 2435 2 2621 1 INV1S $T=825840 477240 1 0 $X=825840 $Y=471820
X922 2651 2 2644 1 INV1S $T=828940 447000 0 180 $X=827700 $Y=441580
X923 2590 2 2660 1 INV1S $T=828320 457080 1 0 $X=828320 $Y=451660
X924 2626 2 2662 1 INV1S $T=830800 416760 1 0 $X=830800 $Y=411340
X925 2661 2 2657 1 INV1S $T=832040 447000 0 180 $X=830800 $Y=441580
X926 2613 2 2667 1 INV1S $T=831420 426840 0 0 $X=831420 $Y=426460
X927 2635 2 2669 1 INV1S $T=832660 426840 1 0 $X=832660 $Y=421420
X928 2619 2 2674 1 INV1S $T=833900 426840 1 0 $X=833900 $Y=421420
X929 2617 2 2676 1 INV1S $T=834520 416760 1 0 $X=834520 $Y=411340
X930 2566 2 2677 1 INV1S $T=834520 457080 1 0 $X=834520 $Y=451660
X931 359 2 2716 1 INV1S $T=843820 537720 0 0 $X=843820 $Y=537340
X932 2693 2 2714 1 INV1S $T=845060 517560 0 0 $X=845060 $Y=517180
X933 2703 2 2719 1 INV1S $T=845060 527640 0 0 $X=845060 $Y=527260
X934 2724 2 2725 1 INV1S $T=847540 517560 0 0 $X=847540 $Y=517180
X935 2700 2 2738 1 INV1S $T=849400 517560 0 0 $X=849400 $Y=517180
X936 2733 2 2752 1 INV1S $T=853740 487320 1 0 $X=853740 $Y=481900
X937 2750 2 2756 1 INV1S $T=858700 497400 1 0 $X=858700 $Y=491980
X938 2758 2 2771 1 INV1S $T=861800 497400 0 0 $X=861800 $Y=497020
X939 2759 2 2767 1 INV1S $T=861800 507480 0 0 $X=861800 $Y=507100
X940 2751 2 2794 1 INV1S $T=866140 487320 0 0 $X=866140 $Y=486940
X941 2778 2 2781 1 INV1S $T=867380 507480 1 0 $X=867380 $Y=502060
X942 371 2 379 1 INV1S $T=868620 537720 0 0 $X=868620 $Y=537340
X943 2773 2 2793 1 INV1S $T=869240 517560 1 0 $X=869240 $Y=512140
X944 378 2 385 1 INV1S $T=876680 527640 0 0 $X=876680 $Y=527260
X945 2817 2 2824 1 INV1S $T=877920 487320 0 0 $X=877920 $Y=486940
X946 2809 2 2835 1 INV1S $T=879160 517560 0 0 $X=879160 $Y=517180
X947 386 2 2846 1 INV1S $T=879160 537720 0 0 $X=879160 $Y=537340
X948 2834 2 2842 1 INV1S $T=881640 487320 0 0 $X=881640 $Y=486940
X949 381 2 2854 1 INV1S $T=881640 537720 1 0 $X=881640 $Y=532300
X950 2799 2 2861 1 INV1S $T=882880 497400 1 0 $X=882880 $Y=491980
X951 2825 2 2848 1 INV1S $T=882880 507480 1 0 $X=882880 $Y=502060
X952 2838 2 2868 1 INV1S $T=889080 507480 1 0 $X=889080 $Y=502060
X953 400 2 2871 1 INV1S $T=891560 396600 0 180 $X=890320 $Y=391180
X954 2806 2 2882 1 INV1S $T=891560 507480 0 0 $X=891560 $Y=507100
X955 398 2 2876 1 INV1S $T=891560 537720 0 0 $X=891560 $Y=537340
X956 407 2 2895 1 INV1S $T=900860 416760 0 180 $X=899620 $Y=411340
X957 2823 2 2920 1 INV1S $T=902720 487320 0 0 $X=902720 $Y=486940
X958 2935 2 2912 1 INV1S $T=907060 517560 1 180 $X=905820 $Y=517180
X959 2902 2 2947 1 INV1S $T=906440 467160 1 0 $X=906440 $Y=461740
X960 2782 2 412 1 INV1S $T=906440 537720 1 0 $X=906440 $Y=532300
X961 2936 2 2939 1 INV1S $T=907060 527640 0 0 $X=907060 $Y=527260
X962 410 2 2949 1 INV1S $T=908920 537720 0 0 $X=908920 $Y=537340
X963 2945 2 2932 1 INV1S $T=910160 517560 1 0 $X=910160 $Y=512140
X964 2929 2 2967 1 INV1S $T=911400 416760 1 0 $X=911400 $Y=411340
X965 2963 2 2942 1 INV1S $T=912640 477240 1 180 $X=911400 $Y=476860
X966 2955 2 2961 1 INV1S $T=911400 527640 1 0 $X=911400 $Y=522220
X967 2948 2 2976 1 INV1S $T=913260 517560 0 0 $X=913260 $Y=517180
X968 2979 2 2982 1 INV1S $T=915740 497400 0 0 $X=915740 $Y=497020
X969 2918 2 2975 1 INV1S $T=916980 527640 1 180 $X=915740 $Y=527260
X970 419 2 2992 1 INV1S $T=916980 507480 1 0 $X=916980 $Y=502060
X971 2965 2 2987 1 INV1S $T=917600 537720 1 0 $X=917600 $Y=532300
X972 2978 2 2996 1 INV1S $T=918220 477240 1 0 $X=918220 $Y=471820
X973 2995 2 3002 1 INV1S $T=918840 537720 1 0 $X=918840 $Y=532300
X974 2997 2 3004 1 INV1S $T=919460 467160 1 0 $X=919460 $Y=461740
X975 3006 2 3000 1 INV1S $T=920700 507480 0 180 $X=919460 $Y=502060
X976 3016 2 3012 1 INV1S $T=925040 517560 0 180 $X=923800 $Y=512140
X977 3017 2 3013 1 INV1S $T=923800 527640 0 0 $X=923800 $Y=527260
X978 3037 2 3011 1 INV1S $T=928140 497400 0 180 $X=926900 $Y=491980
X979 3041 2 3031 1 INV1S $T=929380 507480 0 180 $X=928140 $Y=502060
X980 3027 2 3029 1 INV1S $T=929380 517560 1 0 $X=929380 $Y=512140
X981 405 2 3055 1 INV1S $T=933720 527640 0 0 $X=933720 $Y=527260
X982 3080 2 3078 1 INV1S $T=943640 467160 0 0 $X=943640 $Y=466780
X983 3084 2 3085 1 INV1S $T=946120 457080 0 0 $X=946120 $Y=456700
X984 3087 2 3089 1 INV1S $T=947360 537720 0 0 $X=947360 $Y=537340
X985 3110 2 3144 1 INV1S $T=956660 497400 1 0 $X=956660 $Y=491980
X986 3138 2 3115 1 INV1S $T=959140 467160 0 180 $X=957900 $Y=461740
X987 3150 2 3136 1 INV1S $T=961620 527640 1 180 $X=960380 $Y=527260
X988 3162 2 3135 1 INV1S $T=964100 467160 0 180 $X=962860 $Y=461740
X989 3165 2 3159 1 INV1S $T=966580 467160 1 180 $X=965340 $Y=466780
X990 3187 2 3168 1 INV1S $T=969060 517560 0 180 $X=967820 $Y=512140
X991 3189 2 3185 1 INV1S $T=971540 497400 1 180 $X=970300 $Y=497020
X992 3193 2 3201 1 INV1S $T=981460 497400 0 0 $X=981460 $Y=497020
X993 3206 2 3217 1 INV1S $T=985800 416760 0 0 $X=985800 $Y=416380
X994 3260 2 3234 1 INV1S $T=1006260 426840 1 180 $X=1005020 $Y=426460
X995 3269 2 3245 1 INV1S $T=1007500 447000 1 180 $X=1006260 $Y=446620
X996 3275 2 3252 1 INV1S $T=1012460 416760 1 180 $X=1011220 $Y=416380
X997 3271 2 473 1 INV1S $T=1014940 396600 0 0 $X=1014940 $Y=396220
X998 3277 2 3270 1 INV1S $T=1016180 477240 0 180 $X=1014940 $Y=471820
X999 3278 2 3262 1 INV1S $T=1017420 517560 1 180 $X=1016180 $Y=517180
X1000 3328 2 3318 1 INV1S $T=1038500 406680 0 180 $X=1037260 $Y=401260
X1001 3332 2 3322 1 INV1S $T=1043460 467160 1 180 $X=1042220 $Y=466780
X1002 3340 2 3325 1 INV1S $T=1044080 406680 1 180 $X=1042840 $Y=406300
X1003 3345 2 3314 1 INV1S $T=1048420 467160 1 180 $X=1047180 $Y=466780
X1004 3353 2 3351 1 INV1S $T=1052760 507480 1 180 $X=1051520 $Y=507100
X1005 3370 2 3348 1 INV1S $T=1058340 527640 0 180 $X=1057100 $Y=522220
X1006 3377 2 3358 1 INV1S $T=1060200 507480 0 180 $X=1058960 $Y=502060
X1007 3373 2 3355 1 INV1S $T=1062060 527640 0 180 $X=1060820 $Y=522220
X1008 3378 2 3371 1 INV1S $T=1065160 487320 0 0 $X=1065160 $Y=486940
X1009 3454 2 3466 1 INV1S $T=1111040 416760 0 0 $X=1111040 $Y=416380
X1010 536 539 533 529 2 1 MXL2HS $T=318060 477240 1 180 $X=312480 $Y=476860
X1011 553 548 511 540 2 1 MXL2HS $T=321780 517560 1 180 $X=316200 $Y=517180
X1012 579 569 563 580 2 1 MXL2HS $T=328600 477240 1 0 $X=328600 $Y=471820
X1013 612 615 620 628 2 1 MXL2HS $T=338520 517560 0 0 $X=338520 $Y=517180
X1014 1058 64 1046 994 2 1 MXL2HS $T=440200 537720 1 180 $X=434620 $Y=537340
X1015 69 64 1099 1058 2 1 MXL2HS $T=451980 537720 1 180 $X=446400 $Y=537340
X1016 1222 1132 1213 1169 2 1 MXL2HS $T=476160 416760 0 180 $X=470580 $Y=411340
X1017 1230 1132 1217 1076 2 1 MXL2HS $T=478640 416760 1 180 $X=473060 $Y=416380
X1018 1257 1233 1246 1173 2 1 MXL2HS $T=485460 416760 1 180 $X=479880 $Y=416380
X1019 1261 1233 1259 1120 2 1 MXL2HS $T=488560 416760 0 180 $X=482980 $Y=411340
X1020 1268 1233 1252 1261 2 1 MXL2HS $T=490420 436920 0 180 $X=484840 $Y=431500
X1021 1272 1233 1270 1222 2 1 MXL2HS $T=494760 416760 0 180 $X=489180 $Y=411340
X1022 1283 1280 1271 1268 2 1 MXL2HS $T=495380 457080 0 180 $X=489800 $Y=451660
X1023 1284 1233 1277 1230 2 1 MXL2HS $T=496000 416760 1 180 $X=490420 $Y=416380
X1024 1285 1280 1278 1272 2 1 MXL2HS $T=496000 447000 0 180 $X=490420 $Y=441580
X1025 1295 1280 1291 1257 2 1 MXL2HS $T=501580 426840 0 180 $X=496000 $Y=421420
X1026 1301 1280 1281 1284 2 1 MXL2HS $T=503440 436920 1 180 $X=497860 $Y=436540
X1027 99 1297 1288 1294 2 1 MXL2HS $T=504060 537720 0 180 $X=498480 $Y=532300
X1028 94 1297 98 101 2 1 MXL2HS $T=499720 537720 0 0 $X=499720 $Y=537340
X1029 102 1297 1289 1300 2 1 MXL2HS $T=506540 527640 0 180 $X=500960 $Y=522220
X1030 1314 1309 1306 1283 2 1 MXL2HS $T=509020 457080 1 180 $X=503440 $Y=456700
X1031 100 1305 1312 1315 2 1 MXL2HS $T=503440 507480 1 0 $X=503440 $Y=502060
X1032 1320 1280 1311 1295 2 1 MXL2HS $T=510880 436920 1 180 $X=505300 $Y=436540
X1033 1300 1309 1307 1301 2 1 MXL2HS $T=511500 467160 0 180 $X=505920 $Y=461740
X1034 1327 1305 1317 1296 2 1 MXL2HS $T=512740 487320 0 180 $X=507160 $Y=481900
X1035 110 1309 1326 1285 2 1 MXL2HS $T=514600 457080 0 180 $X=509020 $Y=451660
X1036 111 1309 1322 1320 2 1 MXL2HS $T=514600 477240 0 180 $X=509020 $Y=471820
X1037 106 1297 108 111 2 1 MXL2HS $T=509640 537720 0 0 $X=509640 $Y=537340
X1038 107 1297 1324 1314 2 1 MXL2HS $T=510260 527640 1 0 $X=510260 $Y=522220
X1039 1334 1305 1323 1327 2 1 MXL2HS $T=518320 497400 0 180 $X=512740 $Y=491980
X1040 1315 1305 1318 1334 2 1 MXL2HS $T=521420 497400 1 180 $X=515840 $Y=497020
X1041 118 113 1354 125 2 1 MXL2HS $T=533200 527640 1 180 $X=527620 $Y=527260
X1042 119 113 1398 1360 2 1 MXL2HS $T=535060 527640 0 0 $X=535060 $Y=527260
X1043 129 113 1414 137 2 1 MXL2HS $T=535060 537720 0 0 $X=535060 $Y=537340
X1044 126 154 1465 150 2 1 MXL2HS $T=559860 537720 0 180 $X=554280 $Y=532300
X1045 1294 154 1499 165 2 1 MXL2HS $T=565440 537720 0 0 $X=565440 $Y=537340
X1046 1360 154 1555 178 2 1 MXL2HS $T=586520 537720 0 0 $X=586520 $Y=537340
X1047 1741 1735 1751 1662 2 1 MXL2HS $T=620000 416760 1 0 $X=620000 $Y=411340
X1048 1840 1837 1796 197 2 1 MXL2HS $T=647900 527640 0 180 $X=642320 $Y=522220
X1049 1856 1837 1814 199 2 1 MXL2HS $T=651620 537720 0 180 $X=646040 $Y=532300
X1050 1860 206 1829 200 2 1 MXL2HS $T=652860 517560 0 180 $X=647280 $Y=512140
X1051 1861 1837 1824 201 2 1 MXL2HS $T=653480 527640 1 180 $X=647900 $Y=527260
X1052 205 1837 1863 1840 2 1 MXL2HS $T=649760 527640 1 0 $X=649760 $Y=522220
X1053 214 212 1864 1856 2 1 MXL2HS $T=656580 537720 1 180 $X=651000 $Y=537340
X1054 210 206 1877 1860 2 1 MXL2HS $T=652860 517560 1 0 $X=652860 $Y=512140
X1055 219 1837 1878 1861 2 1 MXL2HS $T=659680 527640 1 180 $X=654100 $Y=527260
X1056 1920 206 1912 221 2 1 MXL2HS $T=674560 537720 1 180 $X=668980 $Y=537340
X1057 244 206 1917 1920 2 1 MXL2HS $T=680140 537720 1 180 $X=674560 $Y=537340
X1058 1949 1940 1961 1938 2 1 MXL2HS $T=679520 436920 0 0 $X=679520 $Y=436540
X1059 1947 1940 1962 1967 2 1 MXL2HS $T=680140 457080 0 0 $X=680140 $Y=456700
X1060 2246 2267 2293 2242 2 1 MXL2HS $T=744000 406680 0 0 $X=744000 $Y=406300
X1061 2308 2254 2284 2245 2 1 MXL2HS $T=749580 467160 0 180 $X=744000 $Y=461740
X1062 3322 480 3317 3314 2 1 MXL2HS $T=1038500 467160 1 180 $X=1032920 $Y=466780
X1063 3318 480 3305 3325 2 1 MXL2HS $T=1035400 406680 0 0 $X=1035400 $Y=406300
X1064 3348 483 3309 3355 2 1 MXL2HS $T=1049040 527640 1 0 $X=1049040 $Y=522220
X1065 3351 483 3266 3358 2 1 MXL2HS $T=1050280 507480 1 0 $X=1050280 $Y=502060
X1066 3454 3419 1 2 INV8 $T=1111660 426840 1 180 $X=1105460 $Y=426460
X1067 141 61 1 2 INV12CK $T=542500 517560 0 180 $X=532580 $Y=512140
X1068 2535 204 1 2 INV12CK $T=802900 487320 0 180 $X=792980 $Y=481900
X1069 2535 344 1 2 INV12CK $T=834520 487320 0 180 $X=824600 $Y=481900
X1070 2535 232 1 2 INV12CK $T=833900 537720 0 0 $X=833900 $Y=537340
X1071 364 2535 1 2 INV12CK $T=847540 537720 0 0 $X=847540 $Y=537340
X1072 425 2813 1 2 INV12CK $T=934340 426840 1 180 $X=924420 $Y=426460
X1073 424 3028 1 2 INV12CK $T=925040 447000 0 0 $X=925040 $Y=446620
X1074 3028 425 1 2 INV12CK $T=925660 416760 0 0 $X=925660 $Y=416380
X1075 3028 453 1 2 INV12CK $T=982080 406680 0 0 $X=982080 $Y=406300
X1076 3028 3241 1 2 INV12CK $T=995100 426840 0 0 $X=995100 $Y=426460
X1077 3241 3151 1 2 INV12CK $T=1018660 426840 1 180 $X=1008740 $Y=426460
X1078 3241 3327 1 2 INV12CK $T=1045940 436920 0 0 $X=1045940 $Y=436540
X1079 3241 485 1 2 INV12CK $T=1058960 426840 0 0 $X=1058960 $Y=426460
X1080 648 623 1 2 523 AN2 $T=347200 507480 0 180 $X=344720 $Y=502060
X1081 672 655 1 2 566 AN2 $T=352780 517560 1 180 $X=350300 $Y=517180
X1082 1088 1074 1 2 1103 AN2 $T=447020 507480 0 0 $X=447020 $Y=507100
X1083 1825 189 1 2 1822 AN2 $T=643560 396600 1 0 $X=643560 $Y=391180
X1084 2050 2066 1 2 2078 AN2 $T=704320 497400 1 0 $X=704320 $Y=491980
X1085 2476 2481 1 2 2491 AN2 $T=787400 426840 0 0 $X=787400 $Y=426460
X1086 361 2716 1 2 2729 AN2 $T=849400 537720 1 0 $X=849400 $Y=532300
X1087 2915 2920 1 2 2921 AN2 $T=903960 507480 1 0 $X=903960 $Y=502060
X1088 3078 3073 1 2 3092 AN2 $T=946120 467160 0 0 $X=946120 $Y=466780
X1089 3115 3086 1 2 3120 AN2 $T=954180 467160 1 0 $X=954180 $Y=461740
X1090 12 512 508 1 2 ND2 $T=301940 537720 1 180 $X=300080 $Y=537340
X1091 519 528 530 1 2 ND2 $T=312480 507480 1 0 $X=312480 $Y=502060
X1092 541 536 538 1 2 ND2 $T=317440 487320 0 180 $X=315580 $Y=481900
X1093 20 551 532 1 2 ND2 $T=321160 537720 1 180 $X=319300 $Y=537340
X1094 560 572 586 1 2 ND2 $T=329840 467160 1 0 $X=329840 $Y=461740
X1095 561 579 588 1 2 ND2 $T=330460 467160 0 0 $X=330460 $Y=466780
X1096 592 538 596 1 2 ND2 $T=332940 487320 1 0 $X=332940 $Y=481900
X1097 599 561 602 1 2 ND2 $T=336040 467160 0 0 $X=336040 $Y=466780
X1098 603 527 600 1 2 ND2 $T=337280 497400 1 0 $X=337280 $Y=491980
X1099 611 560 624 1 2 ND2 $T=339760 457080 0 0 $X=339760 $Y=456700
X1100 617 600 616 1 2 ND2 $T=340380 497400 1 0 $X=340380 $Y=491980
X1101 32 625 31 1 2 ND2 $T=343480 537720 1 180 $X=341620 $Y=537340
X1102 640 634 653 1 2 ND2 $T=345960 447000 0 0 $X=345960 $Y=446620
X1103 652 650 667 1 2 ND2 $T=349680 497400 1 0 $X=349680 $Y=491980
X1104 665 640 670 1 2 ND2 $T=350920 447000 0 0 $X=350920 $Y=446620
X1105 663 623 671 1 2 ND2 $T=354020 507480 1 0 $X=354020 $Y=502060
X1106 697 645 683 1 2 ND2 $T=358980 436920 0 0 $X=358980 $Y=436540
X1107 701 606 700 1 2 ND2 $T=362080 517560 0 0 $X=362080 $Y=517180
X1108 731 738 721 1 2 ND2 $T=367040 436920 0 180 $X=365180 $Y=431500
X1109 752 751 40 1 2 ND2 $T=370760 537720 0 180 $X=368900 $Y=532300
X1110 782 783 756 1 2 ND2 $T=376340 467160 0 180 $X=374480 $Y=461740
X1111 799 742 805 1 2 ND2 $T=381300 426840 0 0 $X=381300 $Y=426460
X1112 838 731 817 1 2 ND2 $T=386880 426840 0 0 $X=386880 $Y=426460
X1113 866 846 839 1 2 ND2 $T=393080 517560 1 0 $X=393080 $Y=512140
X1114 878 900 893 1 2 ND2 $T=397420 426840 0 0 $X=397420 $Y=426460
X1115 880 895 907 1 2 ND2 $T=399280 527640 1 0 $X=399280 $Y=522220
X1116 893 910 896 1 2 ND2 $T=401140 426840 1 0 $X=401140 $Y=421420
X1117 902 907 906 1 2 ND2 $T=403000 527640 1 0 $X=403000 $Y=522220
X1118 878 909 896 1 2 ND2 $T=404860 426840 0 0 $X=404860 $Y=426460
X1119 945 923 954 1 2 ND2 $T=409820 426840 1 0 $X=409820 $Y=421420
X1120 928 954 938 1 2 ND2 $T=414780 426840 1 180 $X=412920 $Y=426460
X1121 958 946 972 1 2 ND2 $T=419120 517560 1 0 $X=419120 $Y=512140
X1122 894 996 848 1 2 ND2 $T=422220 467160 1 180 $X=420360 $Y=466780
X1123 57 983 979 1 2 ND2 $T=422220 406680 0 0 $X=422220 $Y=406300
X1124 967 1002 920 1 2 ND2 $T=426560 507480 0 0 $X=426560 $Y=507100
X1125 60 1011 979 1 2 ND2 $T=430280 406680 0 0 $X=430280 $Y=406300
X1126 1017 1005 1021 1 2 ND2 $T=430280 467160 0 0 $X=430280 $Y=466780
X1127 1027 1013 865 1 2 ND2 $T=431520 497400 1 0 $X=431520 $Y=491980
X1128 57 1062 1055 1 2 ND2 $T=437100 406680 0 0 $X=437100 $Y=406300
X1129 1065 1048 1071 1 2 ND2 $T=440200 457080 0 0 $X=440200 $Y=456700
X1130 4 1064 64 1 2 ND2 $T=441440 527640 1 0 $X=441440 $Y=522220
X1131 1072 1071 1060 1 2 ND2 $T=442680 447000 0 0 $X=442680 $Y=446620
X1132 60 1098 1055 1 2 ND2 $T=444540 406680 0 0 $X=444540 $Y=406300
X1133 811 1109 1077 1 2 ND2 $T=449500 467160 0 180 $X=447640 $Y=461740
X1134 68 1100 979 1 2 ND2 $T=448880 416760 1 0 $X=448880 $Y=411340
X1135 1102 1105 1065 1 2 ND2 $T=449500 457080 1 0 $X=449500 $Y=451660
X1136 74 1136 1132 1 2 ND2 $T=456940 416760 0 180 $X=455080 $Y=411340
X1137 1122 1148 1033 1 2 ND2 $T=458180 436920 1 180 $X=456320 $Y=436540
X1138 1149 1140 1134 1 2 ND2 $T=458180 507480 1 180 $X=456320 $Y=507100
X1139 74 1147 1055 1 2 ND2 $T=458180 416760 1 0 $X=458180 $Y=411340
X1140 1117 1149 1142 1 2 ND2 $T=458800 507480 1 0 $X=458800 $Y=502060
X1141 1003 1163 1155 1 2 ND2 $T=461280 436920 0 180 $X=459420 $Y=431500
X1142 1111 1155 1148 1 2 ND2 $T=459420 436920 0 0 $X=459420 $Y=436540
X1143 1197 1191 1163 1 2 ND2 $T=469340 436920 1 180 $X=467480 $Y=436540
X1144 1171 1198 1186 1 2 ND2 $T=468720 457080 0 0 $X=468720 $Y=456700
X1145 1171 1207 1078 1 2 ND2 $T=473060 457080 1 180 $X=471200 $Y=456700
X1146 1235 1243 1248 1 2 ND2 $T=480500 487320 0 0 $X=480500 $Y=486940
X1147 1247 1248 1239 1 2 ND2 $T=482980 487320 0 180 $X=481120 $Y=481900
X1148 1245 1220 1254 1 2 ND2 $T=482360 457080 1 0 $X=482360 $Y=451660
X1149 1356 1368 1352 1 2 ND2 $T=525760 477240 0 180 $X=523900 $Y=471820
X1150 1368 1363 1353 1 2 ND2 $T=527000 467160 1 180 $X=525140 $Y=466780
X1151 1378 1371 1384 1 2 ND2 $T=530100 426840 1 0 $X=530100 $Y=421420
X1152 128 130 1382 1 2 ND2 $T=533200 396600 0 180 $X=531340 $Y=391180
X1153 1389 1410 1399 1 2 ND2 $T=534440 457080 0 0 $X=534440 $Y=456700
X1154 1374 131 1408 1 2 ND2 $T=535680 447000 0 0 $X=535680 $Y=446620
X1155 1373 1423 1421 1 2 ND2 $T=541260 406680 0 180 $X=539400 $Y=401260
X1156 1483 1490 1474 1 2 ND2 $T=558620 487320 0 180 $X=556760 $Y=481900
X1157 1491 1494 1454 1 2 ND2 $T=561100 487320 1 180 $X=559240 $Y=486940
X1158 1466 1486 1495 1 2 ND2 $T=562340 507480 0 180 $X=560480 $Y=502060
X1159 1482 1504 1450 1 2 ND2 $T=562960 457080 1 180 $X=561100 $Y=456700
X1160 1486 1513 1487 1 2 ND2 $T=561100 497400 1 0 $X=561100 $Y=491980
X1161 1514 161 1519 1 2 ND2 $T=564820 406680 0 0 $X=564820 $Y=406300
X1162 1501 1508 1463 1 2 ND2 $T=564820 487320 0 0 $X=564820 $Y=486940
X1163 1520 1514 1535 1 2 ND2 $T=568540 406680 0 0 $X=568540 $Y=406300
X1164 1537 1559 1533 1 2 ND2 $T=574740 457080 0 180 $X=572880 $Y=451660
X1165 1509 1578 1573 1 2 ND2 $T=579080 507480 1 0 $X=579080 $Y=502060
X1166 1585 1575 1593 1 2 ND2 $T=580320 406680 1 0 $X=580320 $Y=401260
X1167 1512 1579 1580 1 2 ND2 $T=580320 436920 0 0 $X=580320 $Y=436540
X1168 1613 1626 1489 1 2 ND2 $T=588380 416760 0 0 $X=588380 $Y=416380
X1169 1599 1635 1623 1 2 ND2 $T=589000 527640 0 0 $X=589000 $Y=527260
X1170 1642 1657 1646 1 2 ND2 $T=597060 517560 1 180 $X=595200 $Y=517180
X1171 1644 1671 1651 1 2 ND2 $T=599540 527640 1 180 $X=597680 $Y=527260
X1172 1691 1697 1701 1 2 ND2 $T=607600 487320 1 0 $X=607600 $Y=481900
X1173 1702 1711 1558 1 2 ND2 $T=610700 507480 1 180 $X=608840 $Y=507100
X1174 1697 1712 1675 1 2 ND2 $T=610700 487320 0 0 $X=610700 $Y=486940
X1175 1682 1722 1641 1 2 ND2 $T=612560 517560 1 180 $X=610700 $Y=517180
X1176 1688 1738 1680 1 2 ND2 $T=616280 396600 0 0 $X=616280 $Y=396220
X1177 1666 1739 1650 1 2 ND2 $T=616900 487320 1 0 $X=616900 $Y=481900
X1178 1713 1753 1738 1 2 ND2 $T=619380 396600 0 0 $X=619380 $Y=396220
X1179 1634 1754 1650 1 2 ND2 $T=619380 477240 0 0 $X=619380 $Y=476860
X1180 1725 1789 1743 1 2 ND2 $T=631780 507480 0 180 $X=629920 $Y=502060
X1181 1759 1785 1791 1 2 ND2 $T=633640 406680 1 0 $X=633640 $Y=401260
X1182 1742 1806 1670 1 2 ND2 $T=637360 477240 0 180 $X=635500 $Y=471820
X1183 1785 1802 1801 1 2 ND2 $T=639220 406680 0 180 $X=637360 $Y=401260
X1184 1808 1809 1787 1 2 ND2 $T=641700 457080 0 180 $X=639840 $Y=451660
X1185 195 1811 1801 1 2 ND2 $T=642320 396600 1 180 $X=640460 $Y=396220
X1186 1811 1812 1785 1 2 ND2 $T=642320 406680 0 180 $X=640460 $Y=401260
X1187 1841 1859 1847 1 2 ND2 $T=649140 467160 0 0 $X=649140 $Y=466780
X1188 1805 1862 1854 1 2 ND2 $T=651620 426840 1 180 $X=649760 $Y=426460
X1189 1817 1869 1832 1 2 ND2 $T=650380 436920 0 0 $X=650380 $Y=436540
X1190 1889 1921 1927 1 2 ND2 $T=673320 416760 1 0 $X=673320 $Y=411340
X1191 1918 1937 1914 1 2 ND2 $T=678280 426840 0 0 $X=678280 $Y=426460
X1192 1960 1942 1951 1 2 ND2 $T=684480 477240 0 0 $X=684480 $Y=476860
X1193 1969 2010 1988 1 2 ND2 $T=694400 477240 0 180 $X=692540 $Y=471820
X1194 1994 2065 2042 1 2 ND2 $T=703700 457080 1 180 $X=701840 $Y=456700
X1195 2069 2074 269 1 2 ND2 $T=704320 406680 0 0 $X=704320 $Y=406300
X1196 2038 2080 2079 1 2 ND2 $T=704940 416760 0 0 $X=704940 $Y=416380
X1197 2054 2088 2008 1 2 ND2 $T=709280 487320 0 180 $X=707420 $Y=481900
X1198 275 2139 278 1 2 ND2 $T=714240 537720 0 0 $X=714240 $Y=537340
X1199 2145 2124 2120 1 2 ND2 $T=717960 527640 0 180 $X=716100 $Y=522220
X1200 2014 2142 2138 1 2 ND2 $T=718580 457080 1 0 $X=718580 $Y=451660
X1201 1992 2164 2063 1 2 ND2 $T=721060 447000 0 180 $X=719200 $Y=441580
X1202 2157 2165 2124 1 2 ND2 $T=721060 527640 0 180 $X=719200 $Y=522220
X1203 2127 2177 2036 1 2 ND2 $T=722920 527640 1 180 $X=721060 $Y=527260
X1204 281 2179 2152 1 2 ND2 $T=721680 426840 1 0 $X=721680 $Y=421420
X1205 2186 2198 2177 1 2 ND2 $T=728500 527640 1 180 $X=726640 $Y=527260
X1206 2193 2215 2154 1 2 ND2 $T=730360 457080 1 180 $X=728500 $Y=456700
X1207 2110 2205 2116 1 2 ND2 $T=730980 527640 0 180 $X=729120 $Y=522220
X1208 2224 2232 2143 1 2 ND2 $T=734700 517560 1 180 $X=732840 $Y=517180
X1209 1997 2240 2216 1 2 ND2 $T=735940 467160 1 180 $X=734080 $Y=466780
X1210 2216 2262 2169 1 2 ND2 $T=737180 467160 0 0 $X=737180 $Y=466780
X1211 2200 2259 2064 1 2 ND2 $T=740280 517560 1 180 $X=738420 $Y=517180
X1212 2131 2261 2219 1 2 ND2 $T=740900 457080 0 180 $X=739040 $Y=451660
X1213 2270 2275 2261 1 2 ND2 $T=742760 457080 0 180 $X=740900 $Y=451660
X1214 1997 2257 2169 1 2 ND2 $T=740900 467160 1 0 $X=740900 $Y=461740
X1215 2277 2294 2055 1 2 ND2 $T=745860 426840 1 180 $X=744000 $Y=426460
X1216 2109 2299 2286 1 2 ND2 $T=748960 457080 1 180 $X=747100 $Y=456700
X1217 2283 2317 292 1 2 ND2 $T=750200 537720 1 180 $X=748340 $Y=537340
X1218 2296 2318 2183 1 2 ND2 $T=752680 517560 0 180 $X=750820 $Y=512140
X1219 2341 2342 2255 1 2 ND2 $T=755160 517560 0 180 $X=753300 $Y=512140
X1220 296 2375 2356 1 2 ND2 $T=761980 537720 0 180 $X=760120 $Y=532300
X1221 2373 2381 2328 1 2 ND2 $T=763840 507480 1 180 $X=761980 $Y=507100
X1222 2378 2383 2363 1 2 ND2 $T=764460 447000 0 180 $X=762600 $Y=441580
X1223 2307 299 297 1 2 ND2 $T=765080 396600 0 180 $X=763220 $Y=391180
X1224 2347 2384 2353 1 2 ND2 $T=766320 457080 1 180 $X=764460 $Y=456700
X1225 2354 2382 2384 1 2 ND2 $T=764460 467160 0 0 $X=764460 $Y=466780
X1226 300 2403 301 1 2 ND2 $T=770040 537720 1 180 $X=768180 $Y=537340
X1227 2393 2417 2339 1 2 ND2 $T=773760 507480 0 180 $X=771900 $Y=502060
X1228 2391 2422 2401 1 2 ND2 $T=773760 517560 0 180 $X=771900 $Y=512140
X1229 299 2436 2419 1 2 ND2 $T=776860 396600 0 180 $X=775000 $Y=391180
X1230 2416 2470 2456 1 2 ND2 $T=783060 436920 1 180 $X=781200 $Y=436540
X1231 2443 2476 2379 1 2 ND2 $T=783060 416760 0 0 $X=783060 $Y=416380
X1232 2432 2477 2429 1 2 ND2 $T=786160 426840 0 180 $X=784300 $Y=421420
X1233 2456 2473 2477 1 2 ND2 $T=784920 447000 1 0 $X=784920 $Y=441580
X1234 2418 2497 2471 1 2 ND2 $T=788020 537720 0 180 $X=786160 $Y=532300
X1235 2471 2485 313 1 2 ND2 $T=786780 527640 0 0 $X=786780 $Y=527260
X1236 312 2495 2496 1 2 ND2 $T=789880 537720 0 0 $X=789880 $Y=537340
X1237 2502 2517 2396 1 2 ND2 $T=796080 487320 1 180 $X=794220 $Y=486940
X1238 2511 2522 2474 1 2 ND2 $T=797320 477240 0 180 $X=795460 $Y=471820
X1239 2498 2518 2478 1 2 ND2 $T=798560 477240 1 180 $X=796700 $Y=476860
X1240 2504 2540 2490 1 2 ND2 $T=804140 467160 1 180 $X=802280 $Y=466780
X1241 2500 2544 2527 1 2 ND2 $T=807860 457080 0 180 $X=806000 $Y=451660
X1242 2506 2549 2528 1 2 ND2 $T=809100 457080 1 180 $X=807240 $Y=456700
X1243 2547 2554 2526 1 2 ND2 $T=809720 447000 0 180 $X=807860 $Y=441580
X1244 2524 2551 2522 1 2 ND2 $T=809720 477240 1 180 $X=807860 $Y=476860
X1245 2503 2570 2529 1 2 ND2 $T=812820 467160 0 180 $X=810960 $Y=461740
X1246 2543 2567 2574 1 2 ND2 $T=811580 436920 0 0 $X=811580 $Y=436540
X1247 2572 2586 2525 1 2 ND2 $T=815920 426840 0 180 $X=814060 $Y=421420
X1248 2578 2601 2580 1 2 ND2 $T=817160 426840 1 180 $X=815300 $Y=426460
X1249 2600 2606 2565 1 2 ND2 $T=819640 457080 0 180 $X=817780 $Y=451660
X1250 2592 2603 2517 1 2 ND2 $T=819640 487320 1 180 $X=817780 $Y=486940
X1251 2605 2602 2570 1 2 ND2 $T=820260 467160 1 180 $X=818400 $Y=466780
X1252 2568 2612 2521 1 2 ND2 $T=820260 477240 0 180 $X=818400 $Y=471820
X1253 2614 2617 2558 1 2 ND2 $T=822120 416760 0 180 $X=820260 $Y=411340
X1254 2604 2610 2563 1 2 ND2 $T=820880 416760 0 0 $X=820880 $Y=416380
X1255 2618 2643 2594 1 2 ND2 $T=827700 406680 0 180 $X=825840 $Y=401260
X1256 2635 2655 2654 1 2 ND2 $T=832660 426840 0 180 $X=830800 $Y=421420
X1257 2587 2666 2567 1 2 ND2 $T=832660 447000 1 0 $X=832660 $Y=441580
X1258 2667 2675 2601 1 2 ND2 $T=835140 426840 1 180 $X=833280 $Y=426460
X1259 2662 2694 2617 1 2 ND2 $T=838860 416760 0 180 $X=837000 $Y=411340
X1260 2701 2703 351 1 2 ND2 $T=839480 527640 1 180 $X=837620 $Y=527260
X1261 2691 2708 2686 1 2 ND2 $T=842580 517560 1 180 $X=840720 $Y=517180
X1262 2715 2724 2723 1 2 ND2 $T=848160 527640 1 0 $X=848160 $Y=522220
X1263 2720 2726 2673 1 2 ND2 $T=851880 497400 1 180 $X=850020 $Y=497020
X1264 2741 2744 2707 1 2 ND2 $T=855600 497400 1 0 $X=855600 $Y=491980
X1265 2758 371 2768 1 2 ND2 $T=861800 527640 0 0 $X=861800 $Y=527260
X1266 2755 2778 2728 1 2 ND2 $T=864900 507480 0 0 $X=864900 $Y=507100
X1267 2779 2786 2748 1 2 ND2 $T=870480 517560 1 180 $X=868620 $Y=517180
X1268 382 381 2764 1 2 ND2 $T=873580 537720 1 180 $X=871720 $Y=537340
X1269 2803 2807 2801 1 2 ND2 $T=874200 517560 1 180 $X=872340 $Y=517180
X1270 2798 2816 2805 1 2 ND2 $T=877300 497400 1 180 $X=875440 $Y=497020
X1271 2815 2812 2800 1 2 ND2 $T=879780 527640 0 180 $X=877920 $Y=522220
X1272 2825 2821 2820 1 2 ND2 $T=879780 507480 1 0 $X=879780 $Y=502060
X1273 2814 2834 2698 1 2 ND2 $T=881020 497400 1 0 $X=881020 $Y=491980
X1274 2856 2855 2761 1 2 ND2 $T=885980 517560 1 180 $X=884120 $Y=517180
X1275 2878 2899 2885 1 2 ND2 $T=894040 487320 0 0 $X=894040 $Y=486940
X1276 410 2916 2924 1 2 ND2 $T=902720 537720 1 0 $X=902720 $Y=532300
X1277 2932 2923 2908 1 2 ND2 $T=905820 517560 0 180 $X=903960 $Y=512140
X1278 2938 2935 2901 1 2 ND2 $T=907680 517560 0 180 $X=905820 $Y=512140
X1279 410 2955 2939 1 2 ND2 $T=908920 527640 0 0 $X=908920 $Y=527260
X1280 2960 2968 2956 1 2 ND2 $T=912640 497400 1 180 $X=910780 $Y=497020
X1281 2987 2936 3001 1 2 ND2 $T=916980 527640 0 0 $X=916980 $Y=527260
X1282 2993 3016 3005 1 2 ND2 $T=923180 517560 0 180 $X=921320 $Y=512140
X1283 2937 2995 415 1 2 ND2 $T=921320 537720 0 0 $X=921320 $Y=537340
X1284 3018 3027 3032 1 2 ND2 $T=923800 517560 0 0 $X=923800 $Y=517180
X1285 3042 3041 3008 1 2 ND2 $T=928760 507480 1 180 $X=926900 $Y=507100
X1286 3085 3090 3049 1 2 ND2 $T=949840 477240 0 180 $X=947980 $Y=471820
X1287 3067 3096 3100 1 2 ND2 $T=949840 467160 0 0 $X=949840 $Y=466780
X1288 437 3122 3111 1 2 ND2 $T=955420 537720 1 180 $X=953560 $Y=537340
X1289 16 513 1 512 2 520 OAI12HS $T=310620 537720 1 180 $X=306900 $Y=537340
X1290 551 25 1 18 2 578 OAI12HS $T=331080 537720 1 180 $X=327360 $Y=537340
X1291 621 629 1 609 2 596 OAI12HS $T=342240 477240 1 180 $X=338520 $Y=476860
X1292 659 645 1 640 2 635 OAI12HS $T=349060 447000 0 180 $X=345340 $Y=441580
X1293 661 658 1 650 2 618 OAI12HS $T=350300 497400 1 180 $X=346580 $Y=497020
X1294 647 606 1 655 2 639 OAI12HS $T=346580 517560 0 0 $X=346580 $Y=517180
X1295 632 642 1 638 2 609 OAI12HS $T=347200 477240 0 0 $X=347200 $Y=476860
X1296 662 25 1 654 2 680 OAI12HS $T=350920 537720 0 0 $X=350920 $Y=537340
X1297 710 711 1 693 2 670 OAI12HS $T=361460 447000 1 180 $X=357740 $Y=446620
X1298 40 37 1 38 2 39 OAI12HS $T=368280 537720 1 180 $X=364560 $Y=537340
X1299 732 715 1 734 2 693 OAI12HS $T=366420 447000 0 0 $X=366420 $Y=446620
X1300 755 754 1 764 2 765 OAI12HS $T=370760 517560 1 0 $X=370760 $Y=512140
X1301 785 769 1 765 2 770 OAI12HS $T=376340 517560 1 180 $X=372620 $Y=517180
X1302 801 766 1 783 2 775 OAI12HS $T=380060 467160 0 180 $X=376340 $Y=461740
X1303 793 44 1 774 2 763 OAI12HS $T=377580 537720 0 0 $X=377580 $Y=537340
X1304 806 756 1 762 2 755 OAI12HS $T=381920 487320 0 180 $X=378200 $Y=481900
X1305 796 794 1 814 2 683 OAI12HS $T=380680 436920 0 0 $X=380680 $Y=436540
X1306 820 44 1 813 2 849 OAI12HS $T=385020 537720 0 0 $X=385020 $Y=537340
X1307 851 826 1 800 2 814 OAI12HS $T=389360 436920 1 180 $X=385640 $Y=436540
X1308 856 844 1 846 2 754 OAI12HS $T=391220 517560 1 180 $X=387500 $Y=517180
X1309 848 852 1 857 2 853 OAI12HS $T=388740 497400 0 0 $X=388740 $Y=497020
X1310 861 868 1 873 2 851 OAI12HS $T=392460 436920 0 0 $X=392460 $Y=436540
X1311 869 891 1 903 2 873 OAI12HS $T=398660 436920 0 0 $X=398660 $Y=436540
X1312 906 902 1 895 2 892 OAI12HS $T=402380 527640 1 180 $X=398660 $Y=527260
X1313 938 928 1 923 2 817 OAI12HS $T=408580 426840 0 180 $X=404860 $Y=421420
X1314 52 979 1 983 2 977 OAI12HS $T=417260 406680 0 0 $X=417260 $Y=406300
X1315 994 53 1 985 2 987 OAI12HS $T=422840 537720 0 180 $X=419120 $Y=532300
X1316 54 979 1 1011 2 1019 OAI12HS $T=425940 406680 0 0 $X=425940 $Y=406300
X1317 63 64 1 1064 2 1068 OAI12HS $T=437720 527640 1 0 $X=437720 $Y=522220
X1318 1076 1055 1 1062 2 1035 OAI12HS $T=443300 406680 1 180 $X=439580 $Y=406300
X1319 67 979 1 1100 2 1094 OAI12HS $T=446400 416760 0 0 $X=446400 $Y=416380
X1320 1120 1055 1 1098 2 1089 OAI12HS $T=451360 406680 1 180 $X=447640 $Y=406300
X1321 1033 1122 1 1084 2 1111 OAI12HS $T=453840 436920 1 180 $X=450120 $Y=436540
X1322 1113 1061 1 1109 2 1108 OAI12HS $T=454460 467160 0 180 $X=450740 $Y=461740
X1323 72 1132 1 1136 2 1144 OAI12HS $T=454460 416760 0 0 $X=454460 $Y=416380
X1324 1169 1165 1 1124 2 1138 OAI12HS $T=463760 416760 0 180 $X=460040 $Y=411340
X1325 1173 1165 1 1147 2 1161 OAI12HS $T=464380 416760 1 180 $X=460660 $Y=416380
X1326 1296 1236 1 1266 2 1279 OAI12HS $T=500340 487320 1 180 $X=496620 $Y=486940
X1327 1446 1451 1 1457 2 1333 OAI12HS $T=548700 426840 1 0 $X=548700 $Y=421420
X1328 1487 1491 1 1513 2 1522 OAI12HS $T=567920 497400 0 180 $X=564200 $Y=491980
X1329 1497 1502 1 1575 2 170 OAI12HS $T=576600 406680 1 0 $X=576600 $Y=401260
X1330 1500 1572 1 1579 2 1551 OAI12HS $T=577220 447000 1 0 $X=577220 $Y=441580
X1331 1587 1549 1 1578 2 1584 OAI12HS $T=582180 507480 1 180 $X=578460 $Y=507100
X1332 175 168 1 177 2 176 OAI12HS $T=587760 396600 1 0 $X=587760 $Y=391180
X1333 1563 1595 1 1635 2 1644 OAI12HS $T=589000 527640 1 0 $X=589000 $Y=522220
X1334 1497 1616 1 1626 2 1663 OAI12HS $T=592100 426840 1 0 $X=592100 $Y=421420
X1335 1661 1588 1 1639 2 1665 OAI12HS $T=602020 467160 0 180 $X=598300 $Y=461740
X1336 1692 1694 1 1665 2 1714 OAI12HS $T=606360 467160 1 0 $X=606360 $Y=461740
X1337 1701 1691 1 1712 2 1706 OAI12HS $T=608840 477240 0 0 $X=608840 $Y=476860
X1338 1680 1688 1 1708 2 1713 OAI12HS $T=613800 396600 1 180 $X=610080 $Y=396220
X1339 1663 1570 1 1720 2 1723 OAI12HS $T=610700 426840 1 0 $X=610700 $Y=421420
X1340 1699 1716 1 1723 2 1735 OAI12HS $T=611320 416760 0 0 $X=611320 $Y=416380
X1341 1528 1592 1 1724 2 1737 OAI12HS $T=611320 457080 1 0 $X=611320 $Y=451660
X1342 1719 1704 1 1711 2 1743 OAI12HS $T=614420 507480 0 0 $X=614420 $Y=507100
X1343 1729 1718 1 1620 2 1779 OAI12HS $T=623720 457080 1 0 $X=623720 $Y=451660
X1344 1700 1757 1 1705 2 1770 OAI12HS $T=624340 436920 0 0 $X=624340 $Y=436540
X1345 1678 1689 1 1746 2 1764 OAI12HS $T=629300 426840 0 180 $X=625580 $Y=421420
X1346 1763 1769 1 1774 2 1791 OAI12HS $T=627440 406680 0 0 $X=627440 $Y=406300
X1347 1662 1735 1 1686 2 1774 OAI12HS $T=628680 416760 1 0 $X=628680 $Y=411340
X1348 1792 1788 1 1779 2 1787 OAI12HS $T=635500 457080 0 180 $X=631780 $Y=451660
X1349 1980 1968 1 2010 2 2011 OAI12HS $T=693160 477240 0 0 $X=693160 $Y=476860
X1350 1971 1990 1 2043 2 2055 OAI12HS $T=696880 426840 0 0 $X=696880 $Y=426460
X1351 2077 2062 1 2074 2 2106 OAI12HS $T=706180 406680 0 0 $X=706180 $Y=406300
X1352 2091 2062 1 2080 2 2118 OAI12HS $T=709280 426840 1 0 $X=709280 $Y=421420
X1353 2104 2119 1 2088 2 2115 OAI12HS $T=714860 487320 0 180 $X=711140 $Y=481900
X1354 2073 2123 1 2124 2 2117 OAI12HS $T=711760 527640 0 0 $X=711760 $Y=527260
X1355 2129 2034 1 2164 2 2181 OAI12HS $T=721680 447000 1 0 $X=721680 $Y=441580
X1356 2228 2217 1 2205 2 2280 OAI12HS $T=737180 527640 1 0 $X=737180 $Y=522220
X1357 2259 2250 1 2232 2 2282 OAI12HS $T=747100 517560 1 180 $X=743380 $Y=517180
X1358 2219 2131 1 2235 2 2270 OAI12HS $T=744000 457080 1 0 $X=744000 $Y=451660
X1359 2288 2244 1 2295 2 2324 OAI12HS $T=745860 436920 0 0 $X=745860 $Y=436540
X1360 2313 2336 1 2299 2 2353 OAI12HS $T=753920 457080 0 0 $X=753920 $Y=456700
X1361 2260 2272 1 2321 2 2358 OAI12HS $T=755160 426840 0 0 $X=755160 $Y=426460
X1362 2273 2348 1 2259 2 2359 OAI12HS $T=755160 527640 1 0 $X=755160 $Y=522220
X1363 2323 2362 1 2324 2 2363 OAI12HS $T=759500 436920 0 0 $X=759500 $Y=436540
X1364 2318 2357 1 2342 2 2364 OAI12HS $T=763220 517560 0 180 $X=759500 $Y=512140
X1365 2370 2361 1 2358 2 2432 OAI12HS $T=762600 426840 0 0 $X=762600 $Y=426460
X1366 2381 2399 1 2417 2 2405 OAI12HS $T=770040 507480 0 0 $X=770040 $Y=507100
X1367 2422 2365 1 2415 2 2435 OAI12HS $T=773760 517560 1 0 $X=773760 $Y=512140
X1368 2387 2441 1 2381 2 2434 OAI12HS $T=778720 507480 1 180 $X=775000 $Y=507100
X1369 2522 2530 1 2540 2 2536 OAI12HS $T=807240 477240 0 180 $X=803520 $Y=471820
X1370 2517 2539 1 2518 2 2542 OAI12HS $T=808480 487320 0 180 $X=804760 $Y=481900
X1371 2505 2573 1 2517 2 2550 OAI12HS $T=814680 487320 1 180 $X=810960 $Y=486940
X1372 2577 2573 1 2545 2 2588 OAI12HS $T=812820 477240 0 0 $X=812820 $Y=476860
X1373 2544 2575 1 2554 2 2579 OAI12HS $T=813440 447000 0 0 $X=813440 $Y=446620
X1374 2570 2582 1 2549 2 2590 OAI12HS $T=813440 457080 0 0 $X=813440 $Y=456700
X1375 2586 2595 1 2610 2 2619 OAI12HS $T=824600 426840 0 180 $X=820880 $Y=421420
X1376 2609 2573 1 2591 2 2622 OAI12HS $T=824600 487320 0 180 $X=820880 $Y=481900
X1377 2606 2571 1 2585 2 2627 OAI12HS $T=821500 457080 1 0 $X=821500 $Y=451660
X1378 2612 2621 1 2571 2 2629 OAI12HS $T=821500 477240 1 0 $X=821500 $Y=471820
X1379 2564 2623 1 2586 2 2598 OAI12HS $T=822120 436920 1 0 $X=822120 $Y=431500
X1380 2617 2625 1 2643 2 2646 OAI12HS $T=825220 416760 1 0 $X=825220 $Y=411340
X1381 2631 2621 1 2632 2 2650 OAI12HS $T=825220 457080 0 0 $X=825220 $Y=456700
X1382 2655 2623 1 2640 2 2648 OAI12HS $T=830180 436920 0 180 $X=826460 $Y=431500
X1383 2613 2640 1 2601 2 2651 OAI12HS $T=827080 426840 0 0 $X=827080 $Y=426460
X1384 2657 2623 1 2644 2 2652 OAI12HS $T=830800 447000 1 180 $X=827080 $Y=446620
X1385 2645 2621 1 2628 2 2663 OAI12HS $T=828940 477240 1 0 $X=828940 $Y=471820
X1386 2566 2660 1 2544 2 2665 OAI12HS $T=830180 457080 1 0 $X=830180 $Y=451660
X1387 2659 2621 1 2668 2 2684 OAI12HS $T=830800 467160 1 0 $X=830800 $Y=461740
X1388 2669 2638 1 2674 2 2690 OAI12HS $T=835760 426840 1 0 $X=835760 $Y=421420
X1389 2658 2638 1 2688 2 2704 OAI12HS $T=838240 416760 0 0 $X=838240 $Y=416380
X1390 2726 2733 1 2744 2 2750 OAI12HS $T=858700 487320 1 180 $X=854980 $Y=486940
X1391 2751 2766 1 2726 2 2762 OAI12HS $T=864280 487320 1 180 $X=860560 $Y=486940
X1392 2771 2766 1 2756 2 2763 OAI12HS $T=864280 497400 0 180 $X=860560 $Y=491980
X1393 2778 2773 1 2786 2 2788 OAI12HS $T=865520 517560 1 0 $X=865520 $Y=512140
X1394 2765 2766 1 2775 2 2796 OAI12HS $T=872960 507480 0 180 $X=869240 $Y=502060
X1395 371 2766 1 378 2 2810 OAI12HS $T=871720 527640 0 0 $X=871720 $Y=527260
X1396 2807 2809 1 2812 2 2818 OAI12HS $T=874820 517560 0 0 $X=874820 $Y=517180
X1397 2834 2799 1 2816 2 2838 OAI12HS $T=882260 497400 0 0 $X=882260 $Y=497020
X1398 2850 376 1 2859 2 393 OAI12HS $T=884120 537720 0 0 $X=884120 $Y=537340
X1399 2806 2868 1 2807 2 2869 OAI12HS $T=890940 507480 1 180 $X=887220 $Y=507100
X1400 2923 2918 1 2913 2 2906 OAI12HS $T=903960 527640 0 180 $X=900240 $Y=522220
X1401 2945 2948 1 2935 2 2933 OAI12HS $T=908300 517560 0 0 $X=908300 $Y=517180
X1402 2951 2970 1 2957 2 2983 OAI12HS $T=912640 477240 1 0 $X=912640 $Y=471820
X1403 2965 420 1 2995 2 2981 OAI12HS $T=916360 537720 0 0 $X=916360 $Y=537340
X1404 2979 3006 1 2968 2 3009 OAI12HS $T=923800 497400 1 180 $X=920080 $Y=497020
X1405 3026 3025 1 3035 2 3043 OAI12HS $T=925040 467160 0 0 $X=925040 $Y=466780
X1406 3116 3045 1 3097 2 3103 OAI12HS $T=953560 487320 1 180 $X=949840 $Y=486940
X1407 3122 3126 1 3132 2 3117 OAI12HS $T=956040 517560 1 0 $X=956040 $Y=512140
X1408 3128 3129 1 3139 2 3121 OAI12HS $T=956660 477240 1 0 $X=956660 $Y=471820
X1409 3109 3119 1 3141 2 3143 OAI12HS $T=956660 537720 1 0 $X=956660 $Y=532300
X1410 3146 3153 1 3156 2 3140 OAI12HS $T=960380 507480 1 0 $X=960380 $Y=502060
X1411 3172 3176 1 3183 2 3166 OAI12HS $T=967820 507480 1 0 $X=967820 $Y=502060
X1412 543 557 1 568 2 NR2T $T=324880 497400 1 0 $X=324880 $Y=491980
X1413 1464 1456 1 1444 2 NR2T $T=553040 467160 1 180 $X=548080 $Y=466780
X1414 1659 1498 1 1640 2 NR2T $T=600780 507480 0 180 $X=595820 $Y=502060
X1415 1765 1698 1 1749 2 NR2T $T=623100 517560 1 0 $X=623100 $Y=512140
X1416 191 1710 1 1753 2 NR2T $T=624960 396600 1 0 $X=624960 $Y=391180
X1417 1776 1725 1 1743 2 NR2T $T=624960 507480 1 0 $X=624960 $Y=502060
X1418 196 191 1 1785 2 NR2T $T=639220 396600 0 180 $X=634260 $Y=391180
X1419 1800 1786 1 1776 2 NR2T $T=639220 507480 0 180 $X=634260 $Y=502060
X1420 1846 1808 1 1787 2 NR2T $T=644180 447000 1 180 $X=639220 $Y=446620
X1421 1857 1846 1 1826 2 NR2T $T=649140 457080 1 180 $X=644180 $Y=456700
X1422 2271 2070 1 2209 2 NR2T $T=739660 416760 0 0 $X=739660 $Y=416380
X1423 2430 2458 1 2450 2 NR2T $T=778100 426840 0 0 $X=778100 $Y=426460
X1424 2458 2449 1 2379 2 NR2T $T=779340 416760 1 0 $X=779340 $Y=411340
X1425 645 1 643 637 2 636 ND3 $T=347200 436920 1 180 $X=344720 $Y=436540
X1426 656 1 633 636 2 613 ND3 $T=349680 436920 0 180 $X=347200 $Y=431500
X1427 910 1 909 799 2 900 ND3 $T=403620 426840 1 180 $X=401140 $Y=426460
X1428 1023 1 811 1086 2 1073 ND3 $T=447640 487320 0 180 $X=445160 $Y=481900
X1429 1112 1 1105 1133 2 1106 ND3 $T=453840 457080 1 0 $X=453840 $Y=451660
X1430 1188 1 1198 1189 2 1207 ND3 $T=468100 457080 1 0 $X=468100 $Y=451660
X1431 1516 1 1538 1561 2 1509 ND3 $T=577840 497400 1 0 $X=577840 $Y=491980
X1432 1739 1 1754 1772 2 1758 ND3 $T=623100 487320 1 0 $X=623100 $Y=481900
X1433 1869 1 1866 1875 2 1828 ND3 $T=653480 436920 0 0 $X=653480 $Y=436540
X1434 2257 1 2262 2264 2 2240 ND3 $T=740280 467160 0 0 $X=740280 $Y=466780
X1435 2456 1 2427 2465 2 2400 ND3 $T=783680 447000 0 180 $X=781200 $Y=441580
X1436 2471 1 2338 2467 2 2448 ND3 $T=785540 537720 0 180 $X=783060 $Y=532300
X1437 2465 1 2477 2487 2 2470 ND3 $T=786780 436920 1 180 $X=784300 $Y=436540
X1438 313 1 2467 2499 2 2497 ND3 $T=789260 537720 1 0 $X=789260 $Y=532300
X1439 518 517 514 2 1 XNR2HS $T=308760 507480 0 180 $X=303180 $Y=502060
X1440 527 525 521 2 1 XNR2HS $T=313720 497400 0 180 $X=308140 $Y=491980
X1441 556 21 23 2 1 XNR2HS $T=321160 537720 0 0 $X=321160 $Y=537340
X1442 544 572 590 2 1 XNR2HS $T=329220 477240 0 0 $X=329220 $Y=476860
X1443 29 578 610 2 1 XNR2HS $T=335420 537720 0 0 $X=335420 $Y=537340
X1444 638 631 602 2 1 XNR2HS $T=345960 467160 1 180 $X=340380 $Y=466780
X1445 632 642 631 2 1 XNR2HS $T=347820 477240 0 180 $X=342240 $Y=471820
X1446 651 646 592 2 1 XNR2HS $T=348440 487320 0 180 $X=342860 $Y=481900
X1447 652 644 616 2 1 XNR2HS $T=348440 497400 0 180 $X=342860 $Y=491980
X1448 634 637 649 2 1 XNR2HS $T=343480 457080 1 0 $X=343480 $Y=451660
X1449 660 657 644 2 1 XNR2HS $T=350920 487320 1 180 $X=345340 $Y=486940
X1450 679 676 646 2 1 XNR2HS $T=355260 487320 0 180 $X=349680 $Y=481900
X1451 625 680 696 2 1 XNR2HS $T=354640 537720 0 0 $X=354640 $Y=537340
X1452 711 706 697 2 1 XNR2HS $T=363320 447000 0 180 $X=357740 $Y=441580
X1453 712 708 698 2 1 XNR2HS $T=363320 507480 0 180 $X=357740 $Y=502060
X1454 707 702 694 2 1 XNR2HS $T=363940 457080 1 180 $X=358360 $Y=456700
X1455 713 714 704 2 1 XNR2HS $T=365180 436920 0 180 $X=359600 $Y=431500
X1456 726 722 632 2 1 XNR2HS $T=367040 487320 0 180 $X=361460 $Y=481900
X1457 710 734 706 2 1 XNR2HS $T=368900 447000 0 180 $X=363320 $Y=441580
X1458 725 736 681 2 1 XNR2HS $T=368900 467160 1 180 $X=363320 $Y=466780
X1459 730 739 708 2 1 XNR2HS $T=369520 507480 0 180 $X=363940 $Y=502060
X1460 728 748 733 2 1 XNR2HS $T=371380 457080 1 180 $X=365800 $Y=456700
X1461 738 684 758 2 1 XNR2HS $T=368280 436920 0 0 $X=368280 $Y=436540
X1462 735 743 748 2 1 XNR2HS $T=374480 467160 0 180 $X=368900 $Y=461740
X1463 772 759 732 2 1 XNR2HS $T=375720 447000 1 180 $X=370140 $Y=446620
X1464 754 755 768 2 1 XNR2HS $T=370140 507480 1 0 $X=370140 $Y=502060
X1465 775 771 734 2 1 XNR2HS $T=376340 447000 0 180 $X=370760 $Y=441580
X1466 717 763 773 2 1 XNR2HS $T=371380 537720 1 0 $X=371380 $Y=532300
X1467 768 764 686 2 1 XNR2HS $T=377580 507480 1 180 $X=372000 $Y=507100
X1468 796 794 779 2 1 XNR2HS $T=380060 436920 1 180 $X=374480 $Y=436540
X1469 800 779 787 2 1 XNR2HS $T=380680 436920 0 180 $X=375100 $Y=431500
X1470 780 803 771 2 1 XNR2HS $T=382540 447000 0 180 $X=376960 $Y=441580
X1471 762 809 750 2 1 XNR2HS $T=383780 477240 1 180 $X=378200 $Y=476860
X1472 762 810 788 2 1 XNR2HS $T=383780 487320 1 180 $X=378200 $Y=486940
X1473 827 821 801 2 1 XNR2HS $T=386260 467160 1 180 $X=380680 $Y=466780
X1474 818 840 800 2 1 XNR2HS $T=389360 447000 0 180 $X=383780 $Y=441580
X1475 812 808 840 2 1 XNR2HS $T=384400 447000 0 0 $X=384400 $Y=446620
X1476 865 809 825 2 1 XNR2HS $T=394320 487320 1 180 $X=388740 $Y=486940
X1477 821 872 822 2 1 XNR2HS $T=396180 477240 0 180 $X=390600 $Y=471820
X1478 804 872 833 2 1 XNR2HS $T=396180 477240 1 180 $X=390600 $Y=476860
X1479 751 849 875 2 1 XNR2HS $T=391220 537720 1 0 $X=391220 $Y=532300
X1480 861 868 881 2 1 XNR2HS $T=392460 436920 1 0 $X=392460 $Y=431500
X1481 903 881 893 2 1 XNR2HS $T=403620 436920 0 180 $X=398040 $Y=431500
X1482 897 916 874 2 1 XNR2HS $T=405480 447000 1 180 $X=399900 $Y=446620
X1483 927 899 776 2 1 XNR2HS $T=407340 497400 0 180 $X=401760 $Y=491980
X1484 927 922 795 2 1 XNR2HS $T=407340 497400 1 180 $X=401760 $Y=497020
X1485 864 920 886 2 1 XNR2HS $T=403620 467160 1 0 $X=403620 $Y=461740
X1486 946 902 883 2 1 XNR2HS $T=411060 527640 0 180 $X=405480 $Y=522220
X1487 958 809 912 2 1 XNR2HS $T=414160 507480 1 180 $X=408580 $Y=507100
X1488 958 810 933 2 1 XNR2HS $T=417260 517560 0 180 $X=411680 $Y=512140
X1489 961 970 679 2 1 XNR2HS $T=417880 487320 1 180 $X=412300 $Y=486940
X1490 938 928 971 2 1 XNR2HS $T=412920 426840 1 0 $X=412920 $Y=421420
X1491 967 804 960 2 1 XNR2HS $T=419120 497400 1 180 $X=413540 $Y=497020
X1492 973 916 935 2 1 XNR2HS $T=419740 457080 1 180 $X=414160 $Y=456700
X1493 973 879 963 2 1 XNR2HS $T=419740 467160 1 180 $X=414160 $Y=466780
X1494 967 922 974 2 1 XNR2HS $T=414780 507480 0 0 $X=414780 $Y=507100
X1495 982 981 836 2 1 XNR2HS $T=420360 527640 0 180 $X=414780 $Y=522220
X1496 973 972 943 2 1 XNR2HS $T=420980 457080 0 180 $X=415400 $Y=451660
X1497 972 897 984 2 1 XNR2HS $T=416020 447000 0 0 $X=416020 $Y=446620
X1498 990 986 970 2 1 XNR2HS $T=423460 487320 1 180 $X=417880 $Y=486940
X1499 973 993 950 2 1 XNR2HS $T=424700 467160 0 180 $X=419120 $Y=461740
X1500 1002 976 982 2 1 XNR2HS $T=426560 507480 1 180 $X=420980 $Y=507100
X1501 967 899 962 2 1 XNR2HS $T=427180 517560 0 180 $X=421600 $Y=512140
X1502 971 945 1003 2 1 XNR2HS $T=422220 426840 1 0 $X=422220 $Y=421420
X1503 995 1009 959 2 1 XNR2HS $T=429660 457080 0 180 $X=424080 $Y=451660
X1504 864 916 1020 2 1 XNR2HS $T=425940 467160 1 0 $X=425940 $Y=461740
X1505 997 1022 1033 2 1 XNR2HS $T=429660 436920 0 0 $X=429660 $Y=436540
X1506 995 1024 1026 2 1 XNR2HS $T=429660 447000 0 0 $X=429660 $Y=446620
X1507 972 864 1040 2 1 XNR2HS $T=432140 467160 1 0 $X=432140 $Y=461740
X1508 1031 1051 1075 2 1 XNR2HS $T=442060 436920 1 0 $X=442060 $Y=431500
X1509 1073 1024 1085 2 1 XNR2HS $T=442060 477240 0 0 $X=442060 $Y=476860
X1510 1065 998 1101 2 1 XNR2HS $T=445160 477240 1 0 $X=445160 $Y=471820
X1511 1095 1009 1113 2 1 XNR2HS $T=448260 467160 0 0 $X=448260 $Y=466780
X1512 1126 1133 1145 2 1 XNR2HS $T=454460 457080 0 0 $X=454460 $Y=456700
X1513 1146 1152 1157 2 1 XNR2HS $T=459420 497400 1 0 $X=459420 $Y=491980
X1514 1145 1158 1171 2 1 XNR2HS $T=460040 457080 0 0 $X=460040 $Y=456700
X1515 1057 1009 1172 2 1 XNR2HS $T=460040 467160 0 0 $X=460040 $Y=466780
X1516 1081 1108 1182 2 1 XNR2HS $T=461900 467160 1 0 $X=461900 $Y=461740
X1517 1168 1175 1185 2 1 XNR2HS $T=462520 517560 1 0 $X=462520 $Y=512140
X1518 1178 1199 1218 2 1 XNR2HS $T=469960 477240 1 0 $X=469960 $Y=471820
X1519 1182 1218 1247 2 1 XNR2HS $T=478020 477240 1 0 $X=478020 $Y=471820
X1520 1262 1269 1274 2 1 XNR2HS $T=487940 487320 0 0 $X=487940 $Y=486940
X1521 1333 1337 1340 2 1 XNR2HS $T=516460 416760 1 0 $X=516460 $Y=411340
X1522 1345 1332 1336 2 1 XNR2HS $T=522040 426840 1 180 $X=516460 $Y=426460
X1523 1349 1340 115 2 1 XNR2HS $T=522660 406680 1 180 $X=517080 $Y=406300
X1524 1336 1329 1342 2 1 XNR2HS $T=517080 426840 1 0 $X=517080 $Y=421420
X1525 1371 1370 1345 2 1 XNR2HS $T=528240 426840 1 180 $X=522660 $Y=426460
X1526 1352 1356 1381 2 1 XNR2HS $T=527620 477240 1 0 $X=527620 $Y=471820
X1527 1374 1388 1359 2 1 XNR2HS $T=534440 447000 1 180 $X=528860 $Y=446620
X1528 1378 1406 1393 2 1 XNR2HS $T=539400 426840 1 180 $X=533820 $Y=426460
X1529 1387 134 1396 2 1 XNR2HS $T=540020 416760 0 180 $X=534440 $Y=411340
X1530 1385 1413 1397 2 1 XNR2HS $T=540020 467160 1 180 $X=534440 $Y=466780
X1531 1401 1374 1412 2 1 XNR2HS $T=537540 436920 0 0 $X=537540 $Y=436540
X1532 1387 1403 1395 2 1 XNR2HS $T=539400 406680 0 0 $X=539400 $Y=406300
X1533 1378 1434 1402 2 1 XNR2HS $T=547460 426840 0 180 $X=541880 $Y=421420
X1534 1378 1436 1376 2 1 XNR2HS $T=548080 426840 1 180 $X=542500 $Y=426460
X1535 1385 1437 1418 2 1 XNR2HS $T=548080 467160 0 180 $X=542500 $Y=461740
X1536 1385 1438 1419 2 1 XNR2HS $T=548080 477240 0 180 $X=542500 $Y=471820
X1537 1387 1439 1448 2 1 XNR2HS $T=545600 406680 0 0 $X=545600 $Y=406300
X1538 1401 1456 1450 2 1 XNR2HS $T=553660 457080 1 180 $X=548080 $Y=456700
X1539 1461 1388 1471 2 1 XNR2HS $T=551180 457080 1 0 $X=551180 $Y=451660
X1540 1437 1456 1473 2 1 XNR2HS $T=551800 467160 1 0 $X=551800 $Y=461740
X1541 1468 1447 155 2 1 XNR2HS $T=553040 396600 1 0 $X=553040 $Y=391180
X1542 131 1453 1468 2 1 XNR2HS $T=554900 396600 0 0 $X=554900 $Y=396220
X1543 1436 1479 1485 2 1 XNR2HS $T=554900 426840 0 0 $X=554900 $Y=426460
X1544 1434 1460 1478 2 1 XNR2HS $T=555520 416760 0 0 $X=555520 $Y=416380
X1545 1384 1460 1489 2 1 XNR2HS $T=555520 436920 1 0 $X=555520 $Y=431500
X1546 1406 1479 1505 2 1 XNR2HS $T=559860 426840 1 0 $X=559860 $Y=421420
X1547 1401 1463 1507 2 1 XNR2HS $T=559860 477240 0 0 $X=559860 $Y=476860
X1548 1436 1500 1512 2 1 XNR2HS $T=561100 436920 0 0 $X=561100 $Y=436540
X1549 1434 1500 1521 2 1 XNR2HS $T=562340 436920 1 0 $X=562340 $Y=431500
X1550 1495 1466 1524 2 1 XNR2HS $T=562340 507480 0 0 $X=562340 $Y=507100
X1551 1516 1388 1530 2 1 XNR2HS $T=564820 467160 1 0 $X=564820 $Y=461740
X1552 1483 134 1533 2 1 XNR2HS $T=565440 447000 0 0 $X=565440 $Y=446620
X1553 1472 1466 1534 2 1 XNR2HS $T=566060 517560 1 0 $X=566060 $Y=512140
X1554 1406 1500 1536 2 1 XNR2HS $T=566680 426840 0 0 $X=566680 $Y=426460
X1555 1493 1531 1540 2 1 XNR2HS $T=567300 477240 1 0 $X=567300 $Y=471820
X1556 1461 1438 1541 2 1 XNR2HS $T=567300 487320 0 0 $X=567300 $Y=486940
X1557 1519 1403 1542 2 1 XNR2HS $T=567920 406680 1 0 $X=567920 $Y=401260
X1558 1519 1411 1546 2 1 XNR2HS $T=569160 436920 0 0 $X=569160 $Y=436540
X1559 1424 1540 1565 2 1 XNR2HS $T=572880 477240 1 0 $X=572880 $Y=471820
X1560 1439 1500 1577 2 1 XNR2HS $T=575360 447000 0 0 $X=575360 $Y=446620
X1561 1556 1495 1560 2 1 XNR2HS $T=575360 517560 1 0 $X=575360 $Y=512140
X1562 1516 1413 1587 2 1 XNR2HS $T=577220 517560 0 0 $X=577220 $Y=517180
X1563 1408 1487 1573 2 1 XNR2HS $T=581560 507480 1 0 $X=581560 $Y=502060
X1564 1427 1586 174 2 1 XNR2HS $T=582180 396600 1 0 $X=582180 $Y=391180
X1565 1457 134 1616 2 1 XNR2HS $T=584040 426840 1 0 $X=584040 $Y=421420
X1566 1638 1361 1662 2 1 XNR2HS $T=595820 416760 0 0 $X=595820 $Y=416380
X1567 1629 1443 1661 2 1 XNR2HS $T=595820 457080 0 0 $X=595820 $Y=456700
X1568 1566 1517 1649 2 1 XNR2HS $T=602020 487320 0 180 $X=596440 $Y=481900
X1569 1631 1518 1676 2 1 XNR2HS $T=598920 497400 0 0 $X=598920 $Y=497020
X1570 1604 1405 1678 2 1 XNR2HS $T=599540 436920 1 0 $X=599540 $Y=431500
X1571 1364 1632 1680 2 1 XNR2HS $T=600160 396600 0 0 $X=600160 $Y=396220
X1572 1668 1591 1682 2 1 XNR2HS $T=600160 517560 0 0 $X=600160 $Y=517180
X1573 1674 1576 1686 2 1 XNR2HS $T=601400 416760 0 0 $X=601400 $Y=416380
X1574 1669 1672 1674 2 1 XNR2HS $T=602640 416760 1 0 $X=602640 $Y=411340
X1575 1430 1628 1700 2 1 XNR2HS $T=605120 436920 0 0 $X=605120 $Y=436540
X1576 1624 1428 1718 2 1 XNR2HS $T=608840 447000 0 0 $X=608840 $Y=446620
X1577 1676 1715 1725 2 1 XNR2HS $T=610700 507480 1 0 $X=610700 $Y=502060
X1578 1650 1634 1726 2 1 XNR2HS $T=611320 487320 1 0 $X=611320 $Y=481900
X1579 1680 1688 1730 2 1 XNR2HS $T=612560 406680 1 0 $X=612560 $Y=401260
X1580 1592 1528 1734 2 1 XNR2HS $T=613180 467160 1 0 $X=613180 $Y=461740
X1581 1342 186 1747 2 1 XNR2HS $T=618760 416760 0 0 $X=618760 $Y=416380
X1582 1708 1730 1759 2 1 XNR2HS $T=622480 406680 1 0 $X=622480 $Y=401260
X1583 1707 1752 1766 2 1 XNR2HS $T=623720 517560 0 0 $X=623720 $Y=517180
X1584 1718 1729 1760 2 1 XNR2HS $T=630540 457080 1 180 $X=624960 $Y=456700
X1585 1620 1760 1771 2 1 XNR2HS $T=624960 467160 0 0 $X=624960 $Y=466780
X1586 1802 195 1813 2 1 XNR2HS $T=637360 406680 0 0 $X=637360 $Y=406300
X1587 1807 1818 1831 2 1 XNR2HS $T=640460 507480 0 0 $X=640460 $Y=507100
X1588 1859 1855 1874 2 1 XNR2HS $T=651000 477240 1 0 $X=651000 $Y=471820
X1589 1865 1868 1876 2 1 XNR2HS $T=652240 457080 0 0 $X=652240 $Y=456700
X1590 1862 1875 1882 2 1 XNR2HS $T=653480 436920 1 0 $X=653480 $Y=431500
X1591 223 224 230 2 1 XNR2HS $T=662780 396600 1 0 $X=662780 $Y=391180
X1592 223 222 1909 2 1 XNR2HS $T=665880 406680 1 0 $X=665880 $Y=401260
X1593 1921 1919 236 2 1 XNR2HS $T=675180 406680 1 180 $X=669600 $Y=406300
X1594 223 1891 1924 2 1 XNR2HS $T=670840 396600 0 0 $X=670840 $Y=396220
X1595 1886 1916 1936 2 1 XNR2HS $T=673940 436920 0 0 $X=673940 $Y=436540
X1596 1943 1960 1969 2 1 XNR2HS $T=681380 487320 1 0 $X=681380 $Y=481900
X1597 1959 1953 1971 2 1 XNR2HS $T=682620 426840 0 0 $X=682620 $Y=426460
X1598 1958 251 1975 2 1 XNR2HS $T=683240 416760 0 0 $X=683240 $Y=416380
X1599 1932 1959 1983 2 1 XNR2HS $T=685100 426840 1 0 $X=685100 $Y=421420
X1600 1966 1953 1984 2 1 XNR2HS $T=685720 457080 0 0 $X=685720 $Y=456700
X1601 1972 1953 1985 2 1 XNR2HS $T=685720 467160 1 0 $X=685720 $Y=461740
X1602 1899 1950 1988 2 1 XNR2HS $T=686340 477240 1 0 $X=686340 $Y=471820
X1603 1972 1916 1980 2 1 XNR2HS $T=692540 477240 1 180 $X=686960 $Y=476860
X1604 1958 1915 2007 2 1 XNR2HS $T=690060 416760 0 0 $X=690060 $Y=416380
X1605 2027 2020 2002 2 1 XNR2HS $T=697500 507480 0 180 $X=691920 $Y=502060
X1606 260 1977 2030 2 1 XNR2HS $T=693780 537720 0 0 $X=693780 $Y=537340
X1607 1958 1897 2047 2 1 XNR2HS $T=696260 416760 0 0 $X=696260 $Y=416380
X1608 2031 1897 2052 2 1 XNR2HS $T=703080 447000 0 0 $X=703080 $Y=446620
X1609 2031 1915 2051 2 1 XNR2HS $T=710520 447000 0 180 $X=704940 $Y=441580
X1610 2031 1898 2077 2 1 XNR2HS $T=705560 416760 1 0 $X=705560 $Y=411340
X1611 2061 1999 2095 2 1 XNR2HS $T=706800 457080 1 0 $X=706800 $Y=451660
X1612 2031 1927 2083 2 1 XNR2HS $T=713620 436920 1 180 $X=708040 $Y=436540
X1613 2033 2095 2109 2 1 XNR2HS $T=708040 457080 0 0 $X=708040 $Y=456700
X1614 273 251 2121 2 1 XNR2HS $T=709900 416760 0 0 $X=709900 $Y=416380
X1615 1994 1915 2129 2 1 XNR2HS $T=711140 436920 1 0 $X=711140 $Y=431500
X1616 273 1898 2146 2 1 XNR2HS $T=714240 416760 1 0 $X=714240 $Y=411340
X1617 2049 2135 2148 2 1 XNR2HS $T=714240 497400 0 0 $X=714240 $Y=497020
X1618 2134 2068 2156 2 1 XNR2HS $T=716100 477240 1 0 $X=716100 $Y=471820
X1619 2016 2082 2185 2 1 XNR2HS $T=721680 477240 1 0 $X=721680 $Y=471820
X1620 1946 2165 2188 2 1 XNR2HS $T=722300 527640 1 0 $X=722300 $Y=522220
X1621 2136 2170 2190 2 1 XNR2HS $T=722920 537720 1 0 $X=722920 $Y=532300
X1622 2156 2185 2199 2 1 XNR2HS $T=724780 477240 0 0 $X=724780 $Y=476860
X1623 2067 2130 2202 2 1 XNR2HS $T=725400 447000 1 0 $X=725400 $Y=441580
X1624 2117 2198 2225 2 1 XNR2HS $T=729740 537720 1 0 $X=729740 $Y=532300
X1625 2203 2202 2235 2 1 XNR2HS $T=732220 447000 0 0 $X=732220 $Y=446620
X1626 2039 2220 2243 2 1 XNR2HS $T=733460 416760 0 0 $X=733460 $Y=416380
X1627 1976 2175 2245 2 1 XNR2HS $T=733460 457080 1 0 $X=733460 $Y=451660
X1628 2001 2207 2251 2 1 XNR2HS $T=734700 396600 0 0 $X=734700 $Y=396220
X1629 2181 2101 2263 2 1 XNR2HS $T=737800 447000 1 0 $X=737800 $Y=441580
X1630 2192 2094 2267 2 1 XNR2HS $T=738420 406680 0 0 $X=738420 $Y=406300
X1631 2210 2055 2288 2 1 XNR2HS $T=742760 436920 1 0 $X=742760 $Y=431500
X1632 2109 2284 2300 2 1 XNR2HS $T=744000 467160 0 0 $X=744000 $Y=466780
X1633 2191 2081 2301 2 1 XNR2HS $T=744620 396600 1 0 $X=744620 $Y=391180
X1634 2278 2289 2304 2 1 XNR2HS $T=744620 497400 1 0 $X=744620 $Y=491980
X1635 2294 2302 2321 2 1 XNR2HS $T=748340 426840 0 0 $X=748340 $Y=426460
X1636 2291 2301 2333 2 1 XNR2HS $T=752680 396600 1 0 $X=752680 $Y=391180
X1637 2295 2330 2346 2 1 XNR2HS $T=752680 447000 1 0 $X=752680 $Y=441580
X1638 2106 2316 2349 2 1 XNR2HS $T=753300 416760 0 0 $X=753300 $Y=416380
X1639 2272 2260 2350 2 1 XNR2HS $T=753920 436920 1 0 $X=753920 $Y=431500
X1640 1995 2213 2352 2 1 XNR2HS $T=754540 406680 1 0 $X=754540 $Y=401260
X1641 294 295 2356 2 1 XNR2HS $T=755160 537720 0 0 $X=755160 $Y=537340
X1642 2306 2359 2388 2 1 XNR2HS $T=761980 527640 1 0 $X=761980 $Y=522220
X1643 2321 2350 2378 2 1 XNR2HS $T=769420 436920 0 180 $X=763840 $Y=431500
X1644 2410 2400 2407 2 1 XNR2HS $T=772520 467160 1 0 $X=772520 $Y=461740
X1645 2423 2421 2442 2 1 XNR2HS $T=774380 527640 0 0 $X=774380 $Y=527260
X1646 2397 2338 2446 2 1 XNR2HS $T=776860 527640 1 0 $X=776860 $Y=522220
X1647 2445 2438 2459 2 1 XNR2HS $T=778100 457080 0 0 $X=778100 $Y=456700
X1648 305 2437 2464 2 1 XNR2HS $T=779340 406680 1 0 $X=779340 $Y=401260
X1649 2408 2412 2472 2 1 XNR2HS $T=781200 517560 0 0 $X=781200 $Y=517180
X1650 2495 2499 2507 2 1 XNR2HS $T=790500 527640 0 0 $X=790500 $Y=527260
X1651 2552 2550 2546 2 1 XNR2HS $T=810340 487320 1 180 $X=804760 $Y=486940
X1652 2557 2588 2608 2 1 XNR2HS $T=816540 477240 0 0 $X=816540 $Y=476860
X1653 2596 2598 2611 2 1 XNR2HS $T=817160 436920 0 0 $X=817160 $Y=436540
X1654 2551 2622 2649 2 1 XNR2HS $T=824600 477240 0 0 $X=824600 $Y=476860
X1655 2602 2629 2672 2 1 XNR2HS $T=830180 477240 0 0 $X=830180 $Y=476860
X1656 2666 2652 2678 2 1 XNR2HS $T=832040 447000 0 0 $X=832040 $Y=446620
X1657 2583 2663 2680 2 1 XNR2HS $T=832660 477240 1 0 $X=832660 $Y=471820
X1658 2675 2648 2683 2 1 XNR2HS $T=833900 436920 1 0 $X=833900 $Y=431500
X1659 2607 2684 2692 2 1 XNR2HS $T=836380 467160 0 0 $X=836380 $Y=466780
X1660 2685 2650 2697 2 1 XNR2HS $T=837000 457080 0 0 $X=837000 $Y=456700
X1661 2694 2690 2710 2 1 XNR2HS $T=839480 426840 1 0 $X=839480 $Y=421420
X1662 2641 2704 2721 2 1 XNR2HS $T=843200 416760 0 0 $X=843200 $Y=416380
X1663 2760 2762 2774 2 1 XNR2HS $T=861180 487320 1 0 $X=861180 $Y=481900
X1664 2776 2763 2787 2 1 XNR2HS $T=864280 497400 1 0 $X=864280 $Y=491980
X1665 2802 2796 2811 2 1 XNR2HS $T=873580 507480 1 0 $X=873580 $Y=502060
X1666 2831 2810 2849 2 1 XNR2HS $T=880400 527640 1 0 $X=880400 $Y=522220
X1667 2826 2858 2878 2 1 XNR2HS $T=887840 487320 0 0 $X=887840 $Y=486940
X1668 2994 2991 2972 2 1 XNR2HS $T=920080 487320 1 180 $X=914500 $Y=486940
X1669 2944 3010 3021 2 1 XNR2HS $T=920700 487320 0 0 $X=920700 $Y=486940
X1670 3036 3053 3054 2 1 XNR2HS $T=934340 507480 0 0 $X=934340 $Y=507100
X1671 1705 1773 1808 1 2 XOR2H $T=634880 447000 1 0 $X=634880 $Y=441580
X1672 2154 2189 2216 1 2 XOR2H $T=724780 467160 0 0 $X=724780 $Y=466780
X1673 508 2 513 12 1 NR2 $T=300080 537720 1 0 $X=300080 $Y=532300
X1674 13 2 516 9 1 NR2 $T=304420 537720 0 0 $X=304420 $Y=537340
X1675 513 2 532 516 1 NR2 $T=311860 537720 0 0 $X=311860 $Y=537340
X1676 575 2 550 585 1 NR2 $T=327980 517560 1 0 $X=327980 $Y=512140
X1677 547 2 570 589 1 NR2 $T=328600 487320 0 0 $X=328600 $Y=486940
X1678 583 2 585 576 1 NR2 $T=331700 517560 1 0 $X=331700 $Y=512140
X1679 27 2 593 551 1 NR2 $T=334180 537720 1 180 $X=332320 $Y=537340
X1680 589 2 587 538 1 NR2 $T=334800 487320 1 180 $X=332940 $Y=486940
X1681 583 2 584 575 1 NR2 $T=332940 517560 0 0 $X=332940 $Y=517180
X1682 592 2 547 596 1 NR2 $T=335420 487320 1 0 $X=335420 $Y=481900
X1683 624 2 574 611 1 NR2 $T=341000 467160 0 180 $X=339140 $Y=461740
X1684 616 2 589 617 1 NR2 $T=339760 487320 0 0 $X=339760 $Y=486940
X1685 618 2 562 622 1 NR2 $T=340380 497400 0 0 $X=340380 $Y=497020
X1686 626 2 630 576 1 NR2 $T=342860 517560 0 180 $X=341000 $Y=512140
X1687 660 2 674 657 1 NR2 $T=353400 487320 0 0 $X=353400 $Y=486940
X1688 683 2 668 697 1 NR2 $T=355880 436920 0 0 $X=355880 $Y=436540
X1689 702 2 687 705 1 NR2 $T=359600 467160 0 0 $X=359600 $Y=466780
X1690 718 2 713 699 1 NR2 $T=364560 426840 1 180 $X=362700 $Y=426460
X1691 725 2 729 741 1 NR2 $T=365800 477240 1 0 $X=365800 $Y=471820
X1692 739 2 727 730 1 NR2 $T=368900 517560 0 180 $X=367040 $Y=512140
X1693 726 2 737 747 1 NR2 $T=367660 487320 1 0 $X=367660 $Y=481900
X1694 745 2 647 740 1 NR2 $T=368900 517560 0 0 $X=368900 $Y=517180
X1695 772 2 728 760 1 NR2 $T=374480 457080 1 180 $X=372620 $Y=456700
X1696 775 2 791 780 1 NR2 $T=376340 447000 0 0 $X=376340 $Y=446620
X1697 817 2 688 838 1 NR2 $T=383780 426840 0 0 $X=383780 $Y=426460
X1698 855 2 803 862 1 NR2 $T=390600 447000 0 0 $X=390600 $Y=446620
X1699 908 2 818 915 1 NR2 $T=402380 447000 1 0 $X=402380 $Y=441580
X1700 914 2 903 919 1 NR2 $T=403620 436920 1 0 $X=403620 $Y=431500
X1701 926 2 862 932 1 NR2 $T=406100 447000 0 0 $X=406100 $Y=446620
X1702 934 2 915 947 1 NR2 $T=407960 436920 0 0 $X=407960 $Y=436540
X1703 943 2 926 936 1 NR2 $T=410440 447000 1 180 $X=408580 $Y=446620
X1704 933 2 930 918 1 NR2 $T=408580 517560 1 0 $X=408580 $Y=512140
X1705 950 2 934 936 1 NR2 $T=411060 447000 0 180 $X=409200 $Y=441580
X1706 950 2 932 956 1 NR2 $T=410440 447000 0 0 $X=410440 $Y=446620
X1707 921 2 939 962 1 NR2 $T=410440 517560 0 0 $X=410440 $Y=517180
X1708 959 2 947 956 1 NR2 $T=412920 436920 1 180 $X=411060 $Y=436540
X1709 936 2 966 959 1 NR2 $T=412920 436920 0 0 $X=412920 $Y=436540
X1710 966 2 919 969 1 NR2 $T=414780 436920 0 0 $X=414780 $Y=436540
X1711 999 2 969 956 1 NR2 $T=424700 447000 0 180 $X=422840 $Y=441580
X1712 1016 2 1008 997 1 NR2 $T=429040 436920 0 180 $X=427180 $Y=431500
X1713 1018 2 986 1023 1 NR2 $T=429040 497400 0 0 $X=429040 $Y=497020
X1714 1012 2 816 1018 1 NR2 $T=430900 507480 0 180 $X=429040 $Y=502060
X1715 1018 2 968 1025 1 NR2 $T=429660 507480 0 0 $X=429660 $Y=507100
X1716 1038 2 807 1018 1 NR2 $T=434620 507480 1 180 $X=432760 $Y=507100
X1717 1029 2 1042 1031 1 NR2 $T=435240 436920 0 0 $X=435240 $Y=436540
X1718 1024 2 1043 975 1 NR2 $T=436480 447000 0 0 $X=436480 $Y=446620
X1719 65 2 1049 790 1 NR2 $T=438340 497400 1 180 $X=436480 $Y=497020
X1720 1051 2 1030 1056 1 NR2 $T=437100 436920 1 0 $X=437100 $Y=431500
X1721 1052 2 1032 1042 1 NR2 $T=437100 436920 0 0 $X=437100 $Y=436540
X1722 1072 2 1066 1060 1 NR2 $T=442060 447000 1 180 $X=440200 $Y=446620
X1723 1024 2 1067 790 1 NR2 $T=442060 497400 1 180 $X=440200 $Y=497020
X1724 1067 2 1074 888 1 NR2 $T=440820 507480 1 0 $X=440820 $Y=502060
X1725 989 2 1091 1023 1 NR2 $T=445160 497400 0 0 $X=445160 $Y=497020
X1726 1038 2 1102 1071 1 NR2 $T=447640 457080 1 0 $X=447640 $Y=451660
X1727 1103 2 1097 1119 1 NR2 $T=450740 517560 1 0 $X=450740 $Y=512140
X1728 1127 2 1126 953 1 NR2 $T=454460 457080 1 180 $X=452600 $Y=456700
X1729 1127 2 1142 1104 1 NR2 $T=458180 487320 0 180 $X=456320 $Y=481900
X1730 1142 2 1130 1117 1 NR2 $T=458180 507480 0 180 $X=456320 $Y=502060
X1731 1081 2 1158 1139 1 NR2 $T=459420 467160 0 180 $X=457560 $Y=461740
X1732 1200 2 1175 1177 1 NR2 $T=466240 507480 1 180 $X=464380 $Y=507100
X1733 1176 2 1200 1151 1 NR2 $T=465000 497400 0 0 $X=465000 $Y=497020
X1734 1146 2 1195 1152 1 NR2 $T=465620 497400 1 0 $X=465620 $Y=491980
X1735 1143 2 1209 1203 1 NR2 $T=473060 406680 0 180 $X=471200 $Y=401260
X1736 1216 2 1208 1210 1 NR2 $T=473680 507480 0 180 $X=471820 $Y=502060
X1737 1199 2 1221 1178 1 NR2 $T=472440 467160 0 0 $X=472440 $Y=466780
X1738 1206 2 1231 1226 1 NR2 $T=475540 447000 0 0 $X=475540 $Y=446620
X1739 1264 2 1269 1263 1 NR2 $T=487940 467160 0 0 $X=487940 $Y=466780
X1740 1333 2 1331 1337 1 NR2 $T=520800 416760 1 180 $X=518940 $Y=416380
X1741 1352 2 1357 1356 1 NR2 $T=526380 477240 1 180 $X=524520 $Y=476860
X1742 1353 2 1328 1372 1 NR2 $T=525760 457080 1 0 $X=525760 $Y=451660
X1743 1413 2 1420 1425 1 NR2 $T=541260 467160 0 0 $X=541260 $Y=466780
X1744 1454 2 135 1425 1 NR2 $T=543740 487320 0 180 $X=541880 $Y=481900
X1745 1472 2 1453 1425 1 NR2 $T=553660 477240 0 180 $X=551800 $Y=471820
X1746 1454 2 1474 1486 1 NR2 $T=554900 487320 0 0 $X=554900 $Y=486940
X1747 1495 2 1491 1466 1 NR2 $T=561100 507480 1 180 $X=559240 $Y=507100
X1748 1425 2 1532 1538 1 NR2 $T=569160 477240 0 0 $X=569160 $Y=476860
X1749 1538 2 1566 1391 1 NR2 $T=574740 477240 1 180 $X=572880 $Y=476860
X1750 1413 2 1596 1583 1 NR2 $T=582800 487320 1 0 $X=582800 $Y=481900
X1751 1602 2 1600 1596 1 NR2 $T=585900 507480 1 180 $X=584040 $Y=507100
X1752 1614 2 1601 1416 1 NR2 $T=586520 467160 0 0 $X=586520 $Y=466780
X1753 1640 2 1646 1560 1 NR2 $T=595820 517560 0 180 $X=593960 $Y=512140
X1754 1644 2 1654 1651 1 NR2 $T=593960 527640 0 0 $X=593960 $Y=527260
X1755 1572 2 1652 1640 1 NR2 $T=596440 517560 1 0 $X=596440 $Y=512140
X1756 1646 2 1664 1642 1 NR2 $T=598300 517560 0 0 $X=598300 $Y=517180
X1757 1624 2 1673 1677 1 NR2 $T=601400 447000 0 0 $X=601400 $Y=446620
X1758 1612 2 1683 1591 1 NR2 $T=602020 517560 1 0 $X=602020 $Y=512140
X1759 1654 2 1685 1679 1 NR2 $T=602020 527640 0 0 $X=602020 $Y=527260
X1760 1671 2 1693 1664 1 NR2 $T=607600 527640 0 180 $X=605740 $Y=522220
X1761 1641 2 1695 1682 1 NR2 $T=608840 517560 1 180 $X=606980 $Y=517180
X1762 1638 2 1696 1660 1 NR2 $T=609460 406680 1 180 $X=607600 $Y=406300
X1763 1703 2 1707 1693 1 NR2 $T=611320 527640 0 180 $X=609460 $Y=522220
X1764 1643 2 1727 1656 1 NR2 $T=615660 497400 1 180 $X=613800 $Y=497020
X1765 174 2 184 179 1 NR2 $T=616900 396600 0 180 $X=615040 $Y=391180
X1766 1706 2 1731 1645 1 NR2 $T=617520 467160 1 180 $X=615660 $Y=466780
X1767 1744 2 1752 1695 1 NR2 $T=622480 517560 1 180 $X=620620 $Y=517180
X1768 1782 2 1790 1765 1 NR2 $T=632400 517560 1 180 $X=630540 $Y=517180
X1769 1791 2 193 1759 1 NR2 $T=635500 396600 1 180 $X=633640 $Y=396220
X1770 1794 2 1815 1783 1 NR2 $T=637980 497400 0 180 $X=636120 $Y=491980
X1771 1786 2 1818 1815 1 NR2 $T=639840 497400 0 0 $X=639840 $Y=497020
X1772 1821 2 1858 1810 1 NR2 $T=648520 487320 0 0 $X=648520 $Y=486940
X1773 1846 2 1865 1873 1 NR2 $T=655340 457080 1 0 $X=655340 $Y=451660
X1774 1900 2 233 1911 1 NR2 $T=668360 416760 0 0 $X=668360 $Y=416380
X1775 1926 2 239 1900 1 NR2 $T=675180 416760 1 180 $X=673320 $Y=416380
X1776 1918 2 1906 1914 1 NR2 $T=674560 426840 0 0 $X=674560 $Y=426460
X1777 1923 2 241 1900 1 NR2 $T=675800 416760 0 0 $X=675800 $Y=416380
X1778 1926 2 1947 1942 1 NR2 $T=677660 457080 0 0 $X=677660 $Y=456700
X1779 1914 2 1938 1933 1 NR2 $T=680140 447000 0 180 $X=678280 $Y=441580
X1780 1948 2 245 1900 1 NR2 $T=680760 416760 1 180 $X=678900 $Y=416380
X1781 1928 2 1949 246 1 NR2 $T=680760 447000 1 0 $X=680760 $Y=441580
X1782 1932 2 1967 1965 1 NR2 $T=681380 467160 1 0 $X=681380 $Y=461740
X1783 1951 2 1957 1960 1 NR2 $T=681380 477240 0 0 $X=681380 $Y=476860
X1784 1924 2 252 237 1 NR2 $T=688200 396600 0 180 $X=686340 $Y=391180
X1785 257 2 1977 1982 1 NR2 $T=690060 537720 1 180 $X=688200 $Y=537340
X1786 1972 2 2004 1954 1 NR2 $T=693780 447000 1 180 $X=691920 $Y=446620
X1787 1983 2 2015 1990 1 NR2 $T=694400 426840 0 180 $X=692540 $Y=421420
X1788 2058 2 2000 2019 1 NR2 $T=697500 497400 0 180 $X=695640 $Y=491980
X1789 1974 2 2059 2047 1 NR2 $T=699980 426840 1 0 $X=699980 $Y=421420
X1790 2057 2 2058 2044 1 NR2 $T=701220 487320 1 0 $X=701220 $Y=481900
X1791 1913 2 268 2042 1 NR2 $T=701840 436920 1 0 $X=701840 $Y=431500
X1792 2066 2 2027 2050 1 NR2 $T=703700 497400 0 180 $X=701840 $Y=491980
X1793 2042 2 2071 1996 1 NR2 $T=704320 467160 0 0 $X=704320 $Y=466780
X1794 2078 2 2045 2027 1 NR2 $T=706180 497400 1 180 $X=704320 $Y=497020
X1795 2072 2 2066 2054 1 NR2 $T=704940 487320 1 0 $X=704940 $Y=481900
X1796 1916 2 2072 2090 1 NR2 $T=706180 477240 0 0 $X=706180 $Y=476860
X1797 2087 2 2099 2096 1 NR2 $T=708040 497400 1 0 $X=708040 $Y=491980
X1798 2104 2 2097 2057 1 NR2 $T=711140 487320 0 180 $X=709280 $Y=481900
X1799 2099 2 2135 2141 1 NR2 $T=714860 497400 1 0 $X=714860 $Y=491980
X1800 2120 2 2123 2145 1 NR2 $T=716720 527640 0 0 $X=716720 $Y=527260
X1801 2093 2 2158 2140 1 NR2 $T=717340 487320 0 0 $X=717340 $Y=486940
X1802 2162 2 2170 2178 1 NR2 $T=722920 537720 0 0 $X=722920 $Y=537340
X1803 2060 2 2184 2021 1 NR2 $T=724780 457080 0 0 $X=724780 $Y=456700
X1804 2187 2 2194 2201 1 NR2 $T=727880 497400 1 0 $X=727880 $Y=491980
X1805 2175 2 2203 2206 1 NR2 $T=728500 457080 1 0 $X=728500 $Y=451660
X1806 2116 2 2217 2110 1 NR2 $T=729740 517560 0 0 $X=729740 $Y=517180
X1807 2207 2 287 2214 1 NR2 $T=731600 396600 1 0 $X=731600 $Y=391180
X1808 2191 2 2248 2081 1 NR2 $T=735320 396600 1 0 $X=735320 $Y=391180
X1809 2143 2 2250 2224 1 NR2 $T=735320 517560 0 0 $X=735320 $Y=517180
X1810 2101 2 2268 2181 1 NR2 $T=737180 436920 0 0 $X=737180 $Y=436540
X1811 2064 2 2273 2200 1 NR2 $T=740900 517560 0 0 $X=740900 $Y=517180
X1812 2276 2 2297 2266 1 NR2 $T=744000 527640 1 180 $X=742140 $Y=527260
X1813 2285 2 2289 2287 1 NR2 $T=746480 487320 0 0 $X=746480 $Y=486940
X1814 2213 2 2291 2292 1 NR2 $T=749580 406680 0 180 $X=747720 $Y=401260
X1815 2183 2 2305 2296 1 NR2 $T=747720 517560 1 0 $X=747720 $Y=512140
X1816 2196 2 2326 2118 1 NR2 $T=751440 426840 1 0 $X=751440 $Y=421420
X1817 2250 2 2334 2273 1 NR2 $T=752680 517560 0 0 $X=752680 $Y=517180
X1818 2322 2 2327 2344 1 NR2 $T=754540 477240 0 0 $X=754540 $Y=476860
X1819 2255 2 2357 2341 1 NR2 $T=756400 517560 1 0 $X=756400 $Y=512140
X1820 296 2 2390 2356 1 NR2 $T=764460 537720 1 0 $X=764460 $Y=532300
X1821 2328 2 2387 2373 1 NR2 $T=765080 507480 0 0 $X=765080 $Y=507100
X1822 2357 2 2391 2305 1 NR2 $T=765080 517560 1 0 $X=765080 $Y=512140
X1823 2243 2 2376 2360 1 NR2 $T=765700 426840 1 0 $X=765700 $Y=421420
X1824 2275 2 2402 2346 1 NR2 $T=767560 457080 0 180 $X=765700 $Y=451660
X1825 2339 2 2399 2393 1 NR2 $T=765700 507480 1 0 $X=765700 $Y=502060
X1826 2399 2 2401 2387 1 NR2 $T=768180 507480 0 0 $X=768180 $Y=507100
X1827 2409 2 2423 2398 1 NR2 $T=773140 537720 0 0 $X=773140 $Y=537340
X1828 2431 2 2445 2380 1 NR2 $T=776240 457080 1 0 $X=776240 $Y=451660
X1829 2387 2 2455 2454 1 NR2 $T=779340 507480 0 0 $X=779340 $Y=507100
X1830 2396 2 2505 2502 1 NR2 $T=790500 487320 0 0 $X=790500 $Y=486940
X1831 2474 2 2512 2511 1 NR2 $T=794840 477240 0 0 $X=794840 $Y=476860
X1832 2490 2 2530 2504 1 NR2 $T=798560 467160 0 0 $X=798560 $Y=466780
X1833 2530 2 2521 2512 1 NR2 $T=802280 477240 0 180 $X=800420 $Y=471820
X1834 2478 2 2539 2498 1 NR2 $T=802900 487320 1 0 $X=802900 $Y=481900
X1835 2529 2 2561 2503 1 NR2 $T=807240 467160 1 0 $X=807240 $Y=461740
X1836 2527 2 2566 2500 1 NR2 $T=809100 457080 1 0 $X=809100 $Y=451660
X1837 2525 2 2564 2572 1 NR2 $T=810340 426840 1 0 $X=810340 $Y=421420
X1838 2528 2 2582 2506 1 NR2 $T=810340 457080 0 0 $X=810340 $Y=456700
X1839 2526 2 2575 2547 1 NR2 $T=810960 447000 1 0 $X=810960 $Y=441580
X1840 2575 2 2565 2566 1 NR2 $T=813440 457080 0 180 $X=811580 $Y=451660
X1841 2539 2 2568 2505 1 NR2 $T=811580 487320 1 0 $X=811580 $Y=481900
X1842 2582 2 2600 2561 1 NR2 $T=817160 467160 1 0 $X=817160 $Y=461740
X1843 2563 2 2595 2604 1 NR2 $T=819020 416760 0 0 $X=819020 $Y=416380
X1844 2580 2 2613 2578 1 NR2 $T=819020 426840 0 0 $X=819020 $Y=426460
X1845 2606 2 2615 2612 1 NR2 $T=819640 457080 1 0 $X=819640 $Y=451660
X1846 2558 2 2626 2614 1 NR2 $T=822740 416760 1 0 $X=822740 $Y=411340
X1847 2594 2 2625 2618 1 NR2 $T=823980 406680 1 0 $X=823980 $Y=401260
X1848 2595 2 2635 2564 1 NR2 $T=824600 426840 1 0 $X=824600 $Y=421420
X1849 2566 2 2647 2637 1 NR2 $T=828320 457080 0 180 $X=826460 $Y=451660
X1850 2625 2 2654 2626 1 NR2 $T=828940 416760 1 0 $X=828940 $Y=411340
X1851 2613 2 2661 2655 1 NR2 $T=830800 436920 1 0 $X=830800 $Y=431500
X1852 2686 2 2693 2691 1 NR2 $T=837620 517560 0 0 $X=837620 $Y=517180
X1853 2707 2 2733 2741 1 NR2 $T=851880 497400 1 0 $X=851880 $Y=491980
X1854 2673 2 2751 2720 1 NR2 $T=853740 497400 0 0 $X=853740 $Y=497020
X1855 2733 2 2758 2751 1 NR2 $T=857460 497400 0 0 $X=857460 $Y=497020
X1856 2728 2 2759 2755 1 NR2 $T=857460 507480 0 0 $X=857460 $Y=507100
X1857 2773 2 2768 2759 1 NR2 $T=863660 517560 0 180 $X=861800 $Y=512140
X1858 2748 2 2773 2779 1 NR2 $T=864280 517560 0 0 $X=864280 $Y=517180
X1859 2805 2 2799 2798 1 NR2 $T=873580 497400 1 180 $X=871720 $Y=497020
X1860 2801 2 2806 2803 1 NR2 $T=874820 517560 0 180 $X=872960 $Y=512140
X1861 2764 2 386 382 1 NR2 $T=876680 537720 1 180 $X=874820 $Y=537340
X1862 2800 2 2809 2815 1 NR2 $T=875440 527640 1 0 $X=875440 $Y=522220
X1863 2809 2 2820 2806 1 NR2 $T=876060 517560 1 0 $X=876060 $Y=512140
X1864 2698 2 2817 2814 1 NR2 $T=877920 497400 1 0 $X=877920 $Y=491980
X1865 2799 2 2825 2817 1 NR2 $T=877920 497400 0 0 $X=877920 $Y=497020
X1866 2806 2 2852 2848 1 NR2 $T=885980 507480 1 180 $X=884120 $Y=507100
X1867 2876 2 2875 2887 1 NR2 $T=890940 537720 1 0 $X=890940 $Y=532300
X1868 2887 2 2873 2856 1 NR2 $T=895280 527640 1 180 $X=893420 $Y=527260
X1869 2885 2 403 2887 1 NR2 $T=894040 537720 1 0 $X=894040 $Y=532300
X1870 2887 2 404 2856 1 NR2 $T=897140 527640 0 180 $X=895280 $Y=522220
X1871 2923 2 2924 2936 1 NR2 $T=904580 527640 0 0 $X=904580 $Y=527260
X1872 2883 2 2970 2942 1 NR2 $T=905820 477240 1 0 $X=905820 $Y=471820
X1873 2901 2 2945 2938 1 NR2 $T=908300 517560 1 0 $X=908300 $Y=512140
X1874 2945 2 2946 2955 1 NR2 $T=909540 527640 1 0 $X=909540 $Y=522220
X1875 2897 2 2951 2947 1 NR2 $T=910160 467160 1 0 $X=910160 $Y=461740
X1876 2965 2 2969 2949 1 NR2 $T=913260 537720 1 180 $X=911400 $Y=537340
X1877 2956 2 2979 2960 1 NR2 $T=913260 497400 0 0 $X=913260 $Y=497020
X1878 415 2 2965 2937 1 NR2 $T=913880 537720 0 0 $X=913880 $Y=537340
X1879 2952 2 3014 2996 1 NR2 $T=920080 477240 1 0 $X=920080 $Y=471820
X1880 2944 2 2999 3009 1 NR2 $T=923180 497400 1 0 $X=923180 $Y=491980
X1881 3025 2 3038 3014 1 NR2 $T=925660 477240 0 180 $X=923800 $Y=471820
X1882 3020 2 3025 3004 1 NR2 $T=926900 467160 0 180 $X=925040 $Y=461740
X1883 3021 2 3050 416 1 NR2 $T=927520 487320 0 0 $X=927520 $Y=486940
X1884 2979 2 3037 3041 1 NR2 $T=928760 497400 0 0 $X=928760 $Y=497020
X1885 3049 2 3088 3085 1 NR2 $T=944880 477240 1 0 $X=944880 $Y=471820
X1886 433 2 3107 3089 1 NR2 $T=949840 537720 0 0 $X=949840 $Y=537340
X1887 3119 2 3111 3107 1 NR2 $T=954800 537720 0 180 $X=952940 $Y=532300
X1888 3065 2 3119 3136 1 NR2 $T=953560 527640 0 0 $X=953560 $Y=527260
X1889 3122 2 3104 3142 1 NR2 $T=956660 507480 0 0 $X=956660 $Y=507100
X1890 3153 2 3130 3127 1 NR2 $T=959140 507480 0 180 $X=957280 $Y=502060
X1891 3098 2 3127 3144 1 NR2 $T=958520 497400 0 0 $X=958520 $Y=497020
X1892 3129 2 3131 3155 1 NR2 $T=960380 477240 0 0 $X=960380 $Y=476860
X1893 3145 2 3155 3135 1 NR2 $T=961000 467160 0 0 $X=961000 $Y=466780
X1894 3148 2 3129 3159 1 NR2 $T=961000 477240 1 0 $X=961000 $Y=471820
X1895 3133 2 3123 3083 1 NR2 $T=963480 426840 0 180 $X=961620 $Y=421420
X1896 3154 2 3137 3112 1 NR2 $T=964720 416760 1 180 $X=962860 $Y=416380
X1897 3157 2 3153 3168 1 NR2 $T=962860 507480 0 0 $X=962860 $Y=507100
X1898 3149 2 3160 3185 1 NR2 $T=964720 497400 0 0 $X=964720 $Y=497020
X1899 3176 2 3147 3160 1 NR2 $T=967200 507480 0 180 $X=965340 $Y=502060
X1900 3191 2 3176 3201 1 NR2 $T=973400 497400 0 0 $X=973400 $Y=497020
X1901 455 2 3222 3215 1 NR2 $T=989520 507480 0 180 $X=987660 $Y=502060
X1902 3221 2 3223 3214 1 NR2 $T=992000 426840 0 180 $X=990140 $Y=421420
X1903 554 2 545 1 546 NR2P $T=319300 467160 0 0 $X=319300 $Y=466780
X1904 565 2 560 1 545 NR2P $T=323640 467160 1 0 $X=323640 $Y=461740
X1905 565 2 574 1 567 NR2P $T=329220 467160 1 180 $X=325500 $Y=466780
X1906 582 2 583 1 558 NR2P $T=328600 507480 0 0 $X=328600 $Y=507100
X1907 595 2 587 1 542 NR2P $T=331700 497400 1 0 $X=331700 $Y=491980
X1908 602 2 599 1 565 NR2P $T=334800 467160 1 0 $X=334800 $Y=461740
X1909 582 2 626 1 598 NR2P $T=340380 507480 1 180 $X=336660 $Y=507100
X1910 639 2 630 1 605 NR2P $T=343480 517560 1 0 $X=343480 $Y=512140
X1911 668 2 659 1 619 NR2P $T=349680 447000 1 0 $X=349680 $Y=441580
X1912 671 2 663 1 607 NR2P $T=350300 507480 1 0 $X=350300 $Y=502060
X1913 670 2 665 1 659 NR2P $T=353400 447000 0 0 $X=353400 $Y=446620
X1914 699 2 688 1 613 NR2P $T=357120 426840 0 0 $X=357120 $Y=426460
X1915 700 2 701 1 583 NR2P $T=357120 517560 0 0 $X=357120 $Y=517180
X1916 787 2 799 1 699 NR2P $T=380060 426840 1 180 $X=376340 $Y=426460
X1917 939 2 930 1 902 NR2P $T=409820 517560 1 180 $X=406100 $Y=517180
X1918 955 2 897 1 1000 NR2P $T=423460 436920 1 0 $X=423460 $Y=431500
X1919 865 2 1027 1 1007 NR2P $T=432760 487320 1 180 $X=429040 $Y=486940
X1920 1030 2 1032 1 928 NR2P $T=430900 436920 1 0 $X=430900 $Y=431500
X1921 1127 2 824 1 1179 NR2P $T=463140 487320 0 180 $X=459420 $Y=481900
X1922 1184 2 1160 1 1165 NR2P $T=463760 406680 1 0 $X=463760 $Y=401260
X1923 1201 2 1180 1 1210 NR2P $T=469960 497400 1 0 $X=469960 $Y=491980
X1924 1181 2 1204 1 1206 NR2P $T=471200 447000 1 0 $X=471200 $Y=441580
X1925 1433 2 1356 1 1445 NR2P $T=548080 477240 1 180 $X=544360 $Y=476860
X1926 1586 2 1569 1 172 NR2P $T=582180 396600 0 180 $X=578460 $Y=391180
X1927 1632 2 1648 1 177 NR2P $T=595200 396600 1 0 $X=595200 $Y=391180
X1928 1604 2 1681 1 1672 NR2P $T=604500 426840 0 180 $X=600780 $Y=421420
X1929 1518 2 1631 1 1675 NR2P $T=605740 497400 0 180 $X=602020 $Y=491980
X1930 1629 2 1690 1 1724 NR2P $T=605740 457080 0 0 $X=605740 $Y=456700
X1931 1628 2 1717 1 1720 NR2P $T=613180 436920 0 180 $X=609460 $Y=431500
X1932 1761 2 1768 1 1786 NR2P $T=629920 497400 0 0 $X=629920 $Y=497020
X1933 1777 2 1799 1 1810 NR2P $T=641080 487320 0 180 $X=637360 $Y=481900
X1934 1714 2 1771 1 1826 NR2P $T=643560 467160 0 180 $X=639840 $Y=461740
X1935 2042 2 1974 1 2060 NR2P $T=698740 447000 0 0 $X=698740 $Y=446620
X1936 2059 2 2015 1 2070 NR2P $T=706180 426840 0 180 $X=702460 $Y=421420
X1937 2134 2 2155 1 2154 NR2P $T=719820 467160 1 180 $X=716100 $Y=466780
X1938 2107 2 2090 1 2125 NR2P $T=716720 467160 1 0 $X=716720 $Y=461740
X1939 2171 2 2182 1 2201 NR2P $T=729120 487320 1 180 $X=725400 $Y=486940
X1940 2220 2 2238 1 2242 NR2P $T=737800 416760 1 0 $X=737800 $Y=411340
X1941 2229 2 288 1 2276 NR2P $T=744000 537720 1 180 $X=740280 $Y=537340
X1942 2208 2 2271 1 2298 NR2P $T=745860 416760 0 180 $X=742140 $Y=411340
X1943 2265 2 2279 1 2285 NR2P $T=745240 477240 0 0 $X=745240 $Y=476860
X1944 2331 2 2343 1 2344 NR2P $T=756400 467160 0 180 $X=752680 $Y=461740
X1945 2307 2 297 1 298 NR2P $T=762600 396600 0 180 $X=758880 $Y=391180
X1946 301 2 300 1 2398 NR2P $T=767560 537720 1 180 $X=763840 $Y=537340
X1947 2363 2 2378 1 2380 NR2P $T=766320 447000 1 0 $X=766320 $Y=441580
X1948 2369 2 2386 1 303 NR2P $T=773140 396600 1 180 $X=769420 $Y=396220
X1949 2402 2 2380 1 2427 NR2P $T=776240 457080 0 180 $X=772520 $Y=451660
X1950 2398 2 2390 1 2448 NR2P $T=778100 537720 0 180 $X=774380 $Y=532300
X1951 2432 2 2429 1 2450 NR2P $T=779340 426840 0 180 $X=775620 $Y=421420
X1952 2724 2 2693 1 2727 NR2P $T=845680 517560 1 0 $X=845680 $Y=512140
X1953 397 2 2866 1 405 NR2P $T=899620 527640 1 180 $X=895900 $Y=527260
X1954 756 761 1 766 743 778 2 MOAI1 $T=371380 467160 0 0 $X=371380 $Y=466780
X1955 756 762 1 767 739 777 2 MOAI1 $T=371380 497400 1 0 $X=371380 $Y=491980
X1956 780 775 1 791 690 797 2 MOAI1 $T=375100 457080 1 0 $X=375100 $Y=451660
X1957 756 795 1 792 695 767 2 MOAI1 $T=380680 497400 0 180 $X=376340 $Y=491980
X1958 815 828 1 837 780 843 2 MOAI1 $T=384400 457080 1 0 $X=384400 $Y=451660
X1959 832 815 1 822 735 843 2 MOAI1 $T=385640 467160 1 0 $X=385640 $Y=461740
X1960 815 819 1 843 685 833 2 MOAI1 $T=385640 477240 1 0 $X=385640 $Y=471820
X1961 834 848 1 823 720 833 2 MOAI1 $T=390600 477240 1 180 $X=386260 $Y=476860
X1962 839 847 1 844 730 860 2 MOAI1 $T=388120 507480 0 0 $X=388120 $Y=507100
X1963 870 863 1 843 812 854 2 MOAI1 $T=394940 457080 0 180 $X=390600 $Y=451660
X1964 877 811 1 886 891 766 2 MOAI1 $T=394940 457080 0 0 $X=394940 $Y=456700
X1965 937 948 1 941 707 935 2 MOAI1 $T=412300 457080 1 180 $X=407960 $Y=456700
X1966 937 929 1 918 703 960 2 MOAI1 $T=407960 497400 0 0 $X=407960 $Y=497020
X1967 937 942 1 941 722 963 2 MOAI1 $T=408580 487320 1 0 $X=408580 $Y=481900
X1968 1021 848 1 1028 1029 1036 2 MOAI1 $T=429660 477240 1 0 $X=429660 $Y=471820
X1969 1116 65 1 1121 1117 1107 2 MOAI1 $T=455700 507480 0 180 $X=451360 $Y=502060
X1970 1059 1115 1 989 1153 1096 2 MOAI1 $T=453840 487320 0 0 $X=453840 $Y=486940
X1971 1079 1057 1 1166 1178 824 2 MOAI1 $T=459420 477240 1 0 $X=459420 $Y=471820
X1972 1183 1079 1 1187 1199 824 2 MOAI1 $T=465000 477240 1 0 $X=465000 $Y=471820
X1973 1079 1141 1 824 1186 1172 2 MOAI1 $T=471820 467160 1 180 $X=467480 $Y=466780
X1974 1394 1373 1 1366 1364 1355 2 MOAI1 $T=529480 396600 1 180 $X=525140 $Y=396220
X1975 1389 1420 1 1375 1424 1425 2 MOAI1 $T=538160 477240 1 0 $X=538160 $Y=471820
X1976 1373 1432 1 1366 1447 1435 2 MOAI1 $T=543740 396600 0 0 $X=543740 $Y=396220
X1977 1373 1429 1 1366 151 1448 2 MOAI1 $T=549320 396600 0 0 $X=549320 $Y=396220
X1978 1451 1473 1 1481 1493 1469 2 MOAI1 $T=555520 477240 1 0 $X=555520 $Y=471820
X1979 1511 1446 1 1497 1496 1484 2 MOAI1 $T=564820 406680 0 180 $X=560480 $Y=401260
X1980 1509 1485 1 1520 163 1527 2 MOAI1 $T=563580 416760 0 0 $X=563580 $Y=416380
X1981 1519 1509 1 1515 162 1520 2 MOAI1 $T=565440 416760 1 0 $X=565440 $Y=411340
X1982 1505 1537 1 1520 164 1510 2 MOAI1 $T=573500 426840 0 180 $X=569160 $Y=421420
X1983 1539 1509 1 1543 1557 1530 2 MOAI1 $T=572260 457080 0 0 $X=572260 $Y=456700
X1984 1509 1554 1 1550 1576 1564 2 MOAI1 $T=582180 416760 1 180 $X=577840 $Y=416380
X1985 1603 1585 1 1615 175 1497 2 MOAI1 $T=584660 406680 1 0 $X=584660 $Y=401260
X1986 1602 1477 1 1572 1630 1633 2 MOAI1 $T=586520 507480 0 0 $X=586520 $Y=507100
X1987 1613 1618 1 1589 1636 1497 2 MOAI1 $T=587140 406680 0 0 $X=587140 $Y=406300
X1988 1625 1613 1 1597 1669 1497 2 MOAI1 $T=588380 416760 1 0 $X=588380 $Y=411340
X1989 1611 1619 1 1637 1650 1572 2 MOAI1 $T=589000 487320 1 0 $X=589000 $Y=481900
X1990 1656 1643 1 1727 1761 1676 2 MOAI1 $T=612560 497400 1 0 $X=612560 $Y=491980
X1991 1645 1706 1 1731 1742 1748 2 MOAI1 $T=615040 477240 1 0 $X=615040 $Y=471820
X1992 1904 1925 1 242 247 1924 2 MOAI1 $T=685100 396600 0 180 $X=680760 $Y=391180
X1993 1925 1939 1 234 1976 1936 2 MOAI1 $T=690060 436920 0 180 $X=685720 $Y=431500
X1994 254 1925 1 242 261 1975 2 MOAI1 $T=688820 396600 1 0 $X=688820 $Y=391180
X1995 1992 1978 1 1996 1997 1984 2 MOAI1 $T=695640 457080 1 180 $X=691300 $Y=456700
X1996 1992 1922 1 1996 2016 2025 2 MOAI1 $T=692540 457080 1 0 $X=692540 $Y=451660
X1997 1986 2029 1 2018 2019 2005 2 MOAI1 $T=698740 487320 1 180 $X=694400 $Y=486940
X1998 2076 2038 1 2083 2101 2062 2 MOAI1 $T=705560 436920 1 0 $X=705560 $Y=431500
X1999 2075 269 1 2089 2094 2062 2 MOAI1 $T=713000 406680 0 180 $X=708660 $Y=401260
X2000 1992 2013 1 2034 2130 2137 2 MOAI1 $T=711760 447000 1 0 $X=711760 $Y=441580
X2001 281 2168 1 2173 2191 282 2 MOAI1 $T=721680 396600 1 0 $X=721680 $Y=391180
X2002 281 2166 1 2034 2192 2146 2 MOAI1 $T=722300 416760 1 0 $X=722300 $Y=411340
X2003 2191 2081 1 2248 290 2274 2 MOAI1 $T=738420 396600 1 0 $X=738420 $Y=391180
X2004 2196 2118 1 2294 2360 2326 2 MOAI1 $T=753920 426840 1 0 $X=753920 $Y=421420
X2005 2873 2811 1 2866 2891 2894 2 MOAI1 $T=892180 497400 0 0 $X=892180 $Y=497020
X2006 2873 3039 1 427 428 3055 2 MOAI1 $T=930620 537720 1 0 $X=930620 $Y=532300
X2007 530 1 534 526 2 ND2P $T=313100 497400 0 0 $X=313100 $Y=497020
X2008 558 1 534 559 2 ND2P $T=323020 507480 0 0 $X=323020 $Y=507100
X2009 577 1 534 591 2 ND2P $T=330460 497400 0 0 $X=330460 $Y=497020
X2010 598 1 534 601 2 ND2P $T=336660 507480 1 180 $X=332940 $Y=507100
X2011 619 1 627 604 2 ND2P $T=341000 447000 1 0 $X=341000 $Y=441580
X2012 618 1 622 519 2 ND2P $T=342240 497400 0 0 $X=342240 $Y=497020
X2013 955 1 897 980 2 ND2P $T=423460 436920 0 180 $X=419740 $Y=431500
X2014 998 1 967 781 2 ND2P $T=423460 507480 1 0 $X=423460 $Y=502060
X2015 1206 1 1197 1227 2 ND2P $T=474920 436920 0 0 $X=474920 $Y=436540
X2016 1245 1 1254 1228 2 ND2P $T=481120 447000 0 0 $X=481120 $Y=446620
X2017 1248 1 1240 1260 2 ND2P $T=484840 487320 1 0 $X=484840 $Y=481900
X2018 1556 1 1572 1595 2 ND2P $T=583420 517560 0 0 $X=583420 $Y=517180
X2019 1753 1 1710 189 2 ND2P $T=624340 396600 0 180 $X=620620 $Y=391180
X2020 1749 1 1698 1756 2 ND2P $T=625580 507480 1 180 $X=621860 $Y=507100
X2021 1793 1 1798 1828 2 ND2P $T=641700 436920 0 180 $X=637980 $Y=431500
X2022 1797 1 1803 1805 2 ND2P $T=642320 426840 0 180 $X=638600 $Y=421420
X2023 1714 1 1771 1841 2 ND2P $T=642320 467160 0 0 $X=642320 $Y=466780
X2024 1810 1 1816 1827 2 ND2P $T=643560 477240 0 0 $X=643560 $Y=476860
X2025 1836 1 1817 1823 2 ND2P $T=645420 436920 0 0 $X=645420 $Y=436540
X2026 1842 1 1800 1838 2 ND2P $T=646660 507480 1 0 $X=646660 $Y=502060
X2027 1800 1 1852 1844 2 ND2P $T=647900 497400 0 0 $X=647900 $Y=497020
X2028 1928 1 1940 1945 2 ND2P $T=677040 447000 0 0 $X=677040 $Y=446620
X2029 2128 1 2142 277 2 ND2P $T=714860 457080 1 0 $X=714860 $Y=451660
X2030 2211 1 2199 2221 2 ND2P $T=734080 487320 0 180 $X=730360 $Y=481900
X2031 2229 1 288 2253 2 ND2P $T=738420 537720 1 180 $X=734700 $Y=537340
X2032 2221 1 2231 2258 2 ND2P $T=740900 487320 1 180 $X=737180 $Y=486940
X2033 2276 1 2283 2314 2 ND2P $T=750820 537720 0 180 $X=747100 $Y=532300
X2034 2344 1 2354 2371 2 ND2P $T=763220 467160 0 180 $X=759500 $Y=461740
X2035 2275 1 2346 2368 2 ND2P $T=765700 457080 0 180 $X=761980 $Y=451660
X2036 2369 1 2386 302 2 ND2P $T=769420 396600 1 180 $X=765700 $Y=396220
X2037 2430 1 2416 2440 2 ND2P $T=775620 436920 0 0 $X=775620 $Y=436540
X2038 2418 1 307 314 2 ND2P $T=789260 537720 1 180 $X=785540 $Y=537340
X2039 685 669 687 1 2 642 MAO222 $T=358360 477240 0 180 $X=353400 $Y=471820
X2040 679 651 676 1 2 617 MAO222 $T=360220 487320 0 180 $X=355260 $Y=481900
X2041 689 686 692 1 2 700 MAO222 $T=363940 517560 0 180 $X=358980 $Y=512140
X2042 735 728 743 1 2 673 MAO222 $T=368900 467160 0 180 $X=363940 $Y=461740
X2043 723 691 737 1 2 657 MAO222 $T=372620 487320 1 180 $X=367660 $Y=486940
X2044 812 808 818 1 2 715 MAO222 $T=384400 447000 1 180 $X=379440 $Y=446620
X2045 986 961 990 1 2 744 MAO222 $T=422220 497400 0 180 $X=417260 $Y=491980
X2046 1453 1447 131 1 2 144 MAO222 $T=551800 396600 0 180 $X=546840 $Y=391180
X2047 1493 1424 1531 1 2 1588 MAO222 $T=576600 467160 0 0 $X=576600 $Y=466780
X2048 1506 1601 1557 1 2 1620 MAO222 $T=582800 467160 1 0 $X=582800 $Y=461740
X2049 1669 1576 1672 1 2 1688 MAO222 $T=600780 406680 0 0 $X=600780 $Y=406300
X2050 2061 1999 2033 1 2 2131 MAO222 $T=709280 447000 0 0 $X=709280 $Y=446620
X2051 2082 2156 2016 1 2 2226 MAO222 $T=728500 477240 1 0 $X=728500 $Y=471820
X2052 2067 2203 2130 1 2 2244 MAO222 $T=731600 447000 1 0 $X=731600 $Y=441580
X2053 2192 2094 2242 1 2 2281 MAO222 $T=738420 406680 1 0 $X=738420 $Y=401260
X2054 611 673 2 681 641 1 599 FA1 $T=342860 467160 1 0 $X=342860 $Y=461740
X2055 665 690 2 694 733 1 624 FA1 $T=368280 457080 0 180 $X=352780 $Y=451660
X2056 638 716 2 720 729 1 676 FA1 $T=353400 477240 0 0 $X=353400 $Y=476860
X2057 622 698 2 724 682 1 663 FA1 $T=353400 497400 0 0 $X=353400 $Y=497020
X2058 652 703 2 695 744 1 682 FA1 $T=370140 497400 0 180 $X=354640 $Y=491980
X2059 701 786 2 789 770 1 745 FA1 $T=365800 527640 1 0 $X=365800 $Y=522220
X2060 660 790 2 781 830 1 724 FA1 $T=387500 497400 1 180 $X=372000 $Y=497020
X2061 689 807 2 798 845 1 789 FA1 $T=391840 517560 0 180 $X=376340 $Y=512140
X2062 712 781 2 816 859 1 764 FA1 $T=393700 507480 0 180 $X=378200 $Y=502060
X2063 740 850 2 853 892 1 831 FA1 $T=379440 527640 0 0 $X=379440 $Y=527260
X2064 850 968 2 906 965 1 981 FA1 $T=405480 527640 0 0 $X=405480 $Y=527260
X2065 945 991 2 992 1008 1 878 FA1 $T=432760 426840 1 180 $X=417260 $Y=426460
X2066 1174 1153 2 1179 1129 1 1239 FA1 $T=464380 487320 1 0 $X=464380 $Y=481900
X2067 140 1383 2 1379 1404 1 1349 FA1 $T=541880 416760 1 180 $X=526380 $Y=416380
X2068 166 1500 2 131 1496 1 157 FA1 $T=575360 396600 0 180 $X=559860 $Y=391180
X2069 158 1551 2 1532 1458 1 171 FA1 $T=563580 396600 0 0 $X=563580 $Y=396220
X2070 1708 1553 2 1636 1696 1 179 FA1 $T=610080 406680 0 180 $X=594580 $Y=401260
X2071 2132 2115 2 2071 2056 1 2211 FA1 $T=714860 487320 1 0 $X=714860 $Y=481900
X2072 2386 2281 2 2251 2333 1 2307 FA1 $T=763840 396600 1 180 $X=748340 $Y=396220
X2073 2449 2337 2 2352 2293 1 2369 FA1 $T=778100 406680 1 180 $X=762600 $Y=406300
X2074 2443 2337 2 2352 2293 1 3490 FA1 $T=778100 416760 0 180 $X=762600 $Y=411340
X2075 546 547 2 1 531 OR2 $T=319920 487320 0 0 $X=319920 $Y=486940
X2076 583 647 2 1 626 OR2 $T=350300 517560 0 180 $X=347820 $Y=512140
X2077 1040 1104 2 1 1106 OR2 $T=448880 457080 0 0 $X=448880 $Y=456700
X2078 1088 1074 2 1 1123 OR2 $T=450740 507480 0 0 $X=450740 $Y=507100
X2079 1090 1065 2 1 1112 OR2 $T=451360 457080 1 0 $X=451360 $Y=451660
X2080 1133 1126 2 1 1164 OR2 $T=458800 457080 1 0 $X=458800 $Y=451660
X2081 1157 1110 2 1 1167 OR2 $T=460040 497400 0 0 $X=460040 $Y=497020
X2082 1162 1189 2 1 1193 OR2 $T=466240 447000 1 0 $X=466240 $Y=441580
X2083 1195 1223 2 1 1229 OR2 $T=474300 497400 1 0 $X=474300 $Y=491980
X2084 1224 1234 2 1 1244 OR2 $T=478020 467160 1 0 $X=478020 $Y=461740
X2085 1247 1239 2 1 1235 OR2 $T=481120 477240 1 180 $X=478640 $Y=476860
X2086 1242 1256 2 1 1245 OR2 $T=482980 457080 0 0 $X=482980 $Y=456700
X2087 1630 1659 2 1 1702 OR2 $T=606360 507480 0 0 $X=606360 $Y=507100
X2088 1775 1772 2 1 1784 OR2 $T=634880 487320 0 180 $X=632400 $Y=481900
X2089 1776 1842 2 1 1853 OR2 $T=646660 507480 0 0 $X=646660 $Y=507100
X2090 1983 1974 2 1 2043 OR2 $T=696260 426840 1 0 $X=696260 $Y=421420
X2091 1913 1916 2 1 2040 OR2 $T=697500 436920 0 0 $X=697500 $Y=436540
X2092 2103 2048 2 1 2126 OR2 $T=711760 497400 1 0 $X=711760 $Y=491980
X2093 2090 2104 2 1 2128 OR2 $T=712380 457080 1 0 $X=712380 $Y=451660
X2094 2132 2158 2 1 2167 OR2 $T=719820 487320 0 0 $X=719820 $Y=486940
X2095 2127 2036 2 1 2186 OR2 $T=723540 527640 0 0 $X=723540 $Y=527260
X2096 2022 2180 2 1 2197 OR2 $T=724780 436920 0 0 $X=724780 $Y=436540
X2097 2543 2574 2 1 2587 OR2 $T=814060 436920 0 0 $X=814060 $Y=436540
X2098 2701 351 2 1 2715 OR2 $T=841340 527640 0 0 $X=841340 $Y=527260
X2099 361 2716 2 1 2723 OR2 $T=845060 537720 0 0 $X=845060 $Y=537340
X2100 397 398 2 1 2865 OR2 $T=890940 537720 1 180 $X=888460 $Y=537340
X2101 2915 2920 2 1 2908 OR2 $T=903340 507480 0 180 $X=900860 $Y=502060
X2102 2926 2910 2 1 3001 OR2 $T=917600 527640 1 0 $X=917600 $Y=522220
X2103 2993 3005 2 1 3008 OR2 $T=919460 507480 0 0 $X=919460 $Y=507100
X2104 3018 3032 2 1 3042 OR2 $T=926280 517560 0 0 $X=926280 $Y=517180
X2105 3078 3073 2 1 3067 OR2 $T=942400 467160 1 180 $X=939920 $Y=466780
X2106 3115 3086 2 1 3100 OR2 $T=952940 467160 0 180 $X=950460 $Y=461740
X2107 3096 3088 2 1 3093 OR2 $T=950460 477240 1 0 $X=950460 $Y=471820
X2108 19 532 2 520 1 18 AOI12HS $T=318680 537720 1 180 $X=314340 $Y=537340
X2109 613 684 2 627 1 675 AOI12HS $T=355260 436920 1 0 $X=355260 $Y=431500
X2110 721 684 2 749 1 714 AOI12HS $T=367040 436920 1 0 $X=367040 $Y=431500
X2111 752 42 2 746 1 774 AOI12HS $T=375720 537720 1 180 $X=371380 $Y=537340
X2112 1009 1007 2 927 1 1036 AOI12HS $T=429040 487320 1 0 $X=429040 $Y=481900
X2113 1168 1167 2 1200 1 1205 AOI12HS $T=466240 507480 1 0 $X=466240 $Y=502060
X2114 1220 1193 2 1206 1 1190 AOI12HS $T=474920 447000 1 180 $X=470580 $Y=446620
X2115 1438 1445 2 1483 1 1481 AOI12HS $T=566060 477240 0 180 $X=561720 $Y=471820
X2116 1833 1784 2 1810 1 1848 AOI12HS $T=644180 487320 0 0 $X=644180 $Y=486940
X2117 1855 1857 2 1817 1 1872 AOI12HS $T=653480 447000 1 180 $X=649140 $Y=446620
X2118 1847 1855 2 1851 1 1868 AOI12HS $T=651000 467160 1 0 $X=651000 $Y=461740
X2119 1953 1938 2 1940 1 1981 AOI12HS $T=683860 447000 1 0 $X=683860 $Y=441580
X2120 2117 2186 2 2212 1 2228 AOI12HS $T=730360 527640 0 0 $X=730360 $Y=527260
X2121 2253 2218 2 2276 1 2312 AOI12HS $T=745240 527640 0 0 $X=745240 $Y=527260
X2122 2280 2334 2 2282 1 2365 AOI12HS $T=759500 517560 1 180 $X=755160 $Y=517180
X2123 2325 2319 2 2344 1 2372 AOI12HS $T=758260 477240 0 0 $X=758260 $Y=476860
X2124 2364 2401 2 2405 1 2415 AOI12HS $T=767560 517560 1 0 $X=767560 $Y=512140
X2125 2389 2338 2 2413 1 2421 AOI12HS $T=770040 527640 0 0 $X=770040 $Y=527260
X2126 2392 2412 2 2406 1 2425 AOI12HS $T=770660 517560 0 0 $X=770660 $Y=517180
X2127 2414 2400 2 2395 1 2438 AOI12HS $T=771900 457080 0 0 $X=771900 $Y=456700
X2128 2338 2448 2 2418 1 2461 AOI12HS $T=778100 537720 1 0 $X=778100 $Y=532300
X2129 2427 2400 2 2416 1 2468 AOI12HS $T=779340 447000 0 0 $X=779340 $Y=446620
X2130 2455 2412 2 2434 1 2475 AOI12HS $T=781200 507480 0 0 $X=781200 $Y=507100
X2131 2391 2412 2 2364 1 2480 AOI12HS $T=781820 517560 1 0 $X=781820 $Y=512140
X2132 2524 2542 2 2534 1 2545 AOI12HS $T=807240 477240 1 180 $X=802900 $Y=476860
X2133 2542 2521 2 2536 1 2571 AOI12HS $T=816540 477240 0 180 $X=812200 $Y=471820
X2134 2590 2565 2 2579 1 2585 AOI12HS $T=817780 457080 0 180 $X=813440 $Y=451660
X2135 2600 2620 2 2590 1 2632 AOI12HS $T=824600 457080 1 180 $X=820260 $Y=456700
X2136 2615 2435 2 2627 1 2623 AOI12HS $T=821500 447000 0 0 $X=821500 $Y=446620
X2137 2615 2435 2 2627 1 2638 AOI12HS $T=822120 447000 1 0 $X=822120 $Y=441580
X2138 2605 2620 2 2597 1 2628 AOI12HS $T=827080 467160 1 180 $X=822740 $Y=466780
X2139 2619 2654 2 2646 1 2640 AOI12HS $T=830800 426840 0 180 $X=826460 $Y=421420
X2140 2587 2651 2 2636 1 2656 AOI12HS $T=830800 436920 1 180 $X=826460 $Y=436540
X2141 2647 2620 2 2665 1 2668 AOI12HS $T=829560 457080 0 0 $X=829560 $Y=456700
X2142 2662 2619 2 2676 1 2688 AOI12HS $T=832040 416760 0 0 $X=832040 $Y=416380
X2143 2729 2715 2 2719 1 2700 AOI12HS $T=850640 527640 1 180 $X=846300 $Y=527260
X2144 2725 2735 2 2738 1 2747 AOI12HS $T=851880 517560 0 0 $X=851880 $Y=517180
X2145 2723 2735 2 2729 1 2742 AOI12HS $T=856220 537720 0 180 $X=851880 $Y=532300
X2146 2767 2750 2 2781 1 2775 AOI12HS $T=863040 507480 1 0 $X=863040 $Y=502060
X2147 373 374 2 375 1 2782 AOI12HS $T=864280 537720 0 0 $X=864280 $Y=537340
X2148 2750 2768 2 2788 1 378 AOI12HS $T=865520 527640 0 0 $X=865520 $Y=527260
X2149 2838 2820 2 2818 1 2839 AOI12HS $T=882880 507480 1 180 $X=878540 $Y=507100
X2150 2824 2858 2 2842 1 2853 AOI12HS $T=887840 487320 1 180 $X=883500 $Y=486940
X2151 2846 385 2 2854 1 2859 AOI12HS $T=883500 537720 1 0 $X=883500 $Y=532300
X2152 2825 2858 2 2838 1 2867 AOI12HS $T=884740 507480 1 0 $X=884740 $Y=502060
X2153 2852 2858 2 2869 1 2864 AOI12HS $T=886600 517560 1 0 $X=886600 $Y=512140
X2154 2908 2912 2 2921 1 2913 AOI12HS $T=899620 517560 1 0 $X=899620 $Y=512140
X2155 2924 408 2 2906 1 2905 AOI12HS $T=903960 527640 1 180 $X=899620 $Y=527260
X2156 2946 412 2 2933 1 2927 AOI12HS $T=908920 527640 0 180 $X=904580 $Y=522220
X2157 410 412 2 408 1 2964 AOI12HS $T=908300 537720 1 0 $X=908300 $Y=532300
X2158 2939 408 2 2975 1 2948 AOI12HS $T=911400 527640 0 0 $X=911400 $Y=527260
X2159 2961 412 2 2976 1 2980 AOI12HS $T=913260 527640 1 0 $X=913260 $Y=522220
X2160 2969 412 2 2981 1 2988 AOI12HS $T=913260 537720 1 0 $X=913260 $Y=532300
X2161 3002 3001 2 3013 1 2918 AOI12HS $T=919460 527640 0 0 $X=919460 $Y=527260
X2162 3031 2992 2 3000 1 2991 AOI12HS $T=926280 507480 0 180 $X=921940 $Y=502060
X2163 3029 3008 2 3012 1 3006 AOI12HS $T=926280 507480 1 180 $X=921940 $Y=507100
X2164 3037 2992 2 3009 1 3010 AOI12HS $T=928140 497400 1 180 $X=923800 $Y=497020
X2165 2983 3038 2 3043 1 3045 AOI12HS $T=926900 477240 1 0 $X=926900 $Y=471820
X2166 3042 2992 2 3029 1 3053 AOI12HS $T=929380 507480 0 0 $X=929380 $Y=507100
X2167 3104 3103 2 3117 1 3094 AOI12HS $T=951700 507480 1 0 $X=951700 $Y=502060
X2168 3092 3100 2 3120 1 3113 AOI12HS $T=952940 467160 0 0 $X=952940 $Y=466780
X2169 3121 3130 2 3140 1 3097 AOI12HS $T=956040 487320 0 0 $X=956040 $Y=486940
X2170 439 3111 2 3143 1 3132 AOI12HS $T=956660 537720 0 0 $X=956660 $Y=537340
X2171 3166 443 2 444 1 3126 AOI12HS $T=965960 517560 0 180 $X=961620 $Y=512140
X2172 528 535 524 2 1 XOR2HS $T=316200 507480 1 180 $X=310620 $Y=507100
X2173 584 571 510 2 1 XOR2HS $T=332320 517560 1 180 $X=326740 $Y=517180
X2174 669 666 641 2 1 XOR2HS $T=352780 467160 1 180 $X=347200 $Y=466780
X2175 678 675 664 2 1 XOR2HS $T=355260 436920 0 180 $X=349680 $Y=431500
X2176 689 686 677 2 1 XOR2HS $T=358360 517560 0 180 $X=352780 $Y=512140
X2177 685 687 666 2 1 XOR2HS $T=358980 467160 1 180 $X=353400 $Y=466780
X2178 692 677 671 2 1 XOR2HS $T=358980 507480 1 180 $X=353400 $Y=507100
X2179 762 784 761 2 1 XOR2HS $T=377580 487320 0 180 $X=372000 $Y=481900
X2180 762 804 782 2 1 XOR2HS $T=382540 477240 0 180 $X=376960 $Y=471820
X2181 836 831 612 2 1 XOR2HS $T=387500 527640 0 180 $X=381920 $Y=522220
X2182 855 862 826 2 1 XOR2HS $T=395560 447000 0 180 $X=389980 $Y=441580
X2183 872 784 834 2 1 XOR2HS $T=395560 487320 0 180 $X=389980 $Y=481900
X2184 47 44 871 2 1 XOR2HS $T=389980 537720 0 0 $X=389980 $Y=537340
X2185 878 876 838 2 1 XOR2HS $T=396800 426840 1 180 $X=391220 $Y=426460
X2186 879 872 832 2 1 XOR2HS $T=396800 467160 0 180 $X=391220 $Y=461740
X2187 883 880 786 2 1 XOR2HS $T=397420 527640 0 180 $X=391840 $Y=522220
X2188 896 893 876 2 1 XOR2HS $T=400520 426840 0 180 $X=394940 $Y=421420
X2189 899 898 887 2 1 XOR2HS $T=401760 497400 0 180 $X=396180 $Y=491980
X2190 901 899 866 2 1 XOR2HS $T=401760 517560 0 180 $X=396180 $Y=512140
X2191 898 809 884 2 1 XOR2HS $T=402380 477240 1 180 $X=396800 $Y=476860
X2192 810 898 889 2 1 XOR2HS $T=402380 487320 1 180 $X=396800 $Y=486940
X2193 864 879 877 2 1 XOR2HS $T=403000 467160 0 180 $X=397420 $Y=461740
X2194 901 810 847 2 1 XOR2HS $T=403000 507480 0 180 $X=397420 $Y=502060
X2195 922 901 867 2 1 XOR2HS $T=406100 517560 1 180 $X=400520 $Y=517180
X2196 908 915 896 2 1 XOR2HS $T=402380 436920 0 0 $X=402380 $Y=436540
X2197 804 898 913 2 1 XOR2HS $T=407960 477240 1 180 $X=402380 $Y=476860
X2198 784 898 911 2 1 XOR2HS $T=407960 487320 0 180 $X=402380 $Y=481900
X2199 898 922 904 2 1 XOR2HS $T=407960 487320 1 180 $X=402380 $Y=486940
X2200 897 920 828 2 1 XOR2HS $T=409200 457080 0 180 $X=403620 $Y=451660
X2201 914 919 940 2 1 XOR2HS $T=405480 436920 1 0 $X=405480 $Y=431500
X2202 958 784 929 2 1 XOR2HS $T=412920 507480 0 180 $X=407340 $Y=502060
X2203 958 821 942 2 1 XOR2HS $T=413540 477240 1 180 $X=407960 $Y=476860
X2204 973 920 948 2 1 XOR2HS $T=417880 467160 0 180 $X=412300 $Y=461740
X2205 952 821 924 2 1 XOR2HS $T=419120 477240 1 180 $X=413540 $Y=476860
X2206 952 879 964 2 1 XOR2HS $T=417880 477240 1 0 $X=417880 $Y=471820
X2207 952 920 1004 2 1 XOR2HS $T=422840 487320 1 0 $X=422840 $Y=481900
X2208 995 998 1001 2 1 XOR2HS $T=429660 447000 1 180 $X=424080 $Y=446620
X2209 1010 916 1044 2 1 XOR2HS $T=432760 487320 0 0 $X=432760 $Y=486940
X2210 993 1057 1021 2 1 XOR2HS $T=441440 467160 1 180 $X=435860 $Y=466780
X2211 1070 993 1077 2 1 XOR2HS $T=440820 467160 1 0 $X=440820 $Y=461740
X2212 1063 1075 1084 2 1 XOR2HS $T=442060 436920 0 0 $X=442060 $Y=436540
X2213 1010 972 1069 2 1 XOR2HS $T=442680 497400 1 0 $X=442680 $Y=491980
X2214 1010 998 1093 2 1 XOR2HS $T=443300 507480 1 0 $X=443300 $Y=502060
X2215 1072 1060 1047 2 1 XOR2HS $T=444540 447000 0 0 $X=444540 $Y=446620
X2216 1010 993 1115 2 1 XOR2HS $T=448260 487320 0 0 $X=448260 $Y=486940
X2217 1009 1010 1116 2 1 XOR2HS $T=448260 497400 1 0 $X=448260 $Y=491980
X2218 1033 1122 1137 2 1 XOR2HS $T=451980 447000 1 0 $X=451980 $Y=441580
X2219 1057 998 1141 2 1 XOR2HS $T=453840 467160 0 0 $X=453840 $Y=466780
X2220 1123 1140 1156 2 1 XOR2HS $T=456320 517560 1 0 $X=456320 $Y=512140
X2221 1084 1137 1162 2 1 XOR2HS $T=457560 447000 1 0 $X=457560 $Y=441580
X2222 1191 1190 1045 2 1 XOR2HS $T=468720 447000 1 180 $X=463140 $Y=446620
X2223 1057 1024 1183 2 1 XOR2HS $T=463140 477240 0 0 $X=463140 $Y=476860
X2224 1186 1078 1214 2 1 XOR2HS $T=468720 467160 1 0 $X=468720 $Y=461740
X2225 1205 1208 1219 2 1 XOR2HS $T=469960 517560 1 0 $X=469960 $Y=512140
X2226 80 1209 85 2 1 XOR2HS $T=472440 396600 1 0 $X=472440 $Y=391180
X2227 1214 1171 1224 2 1 XOR2HS $T=473060 457080 0 0 $X=473060 $Y=456700
X2228 1220 1231 1215 2 1 XOR2HS $T=479260 457080 0 180 $X=473680 $Y=451660
X2229 1240 1243 1237 2 1 XOR2HS $T=483600 497400 0 180 $X=478020 $Y=491980
X2230 1387 1384 1358 2 1 XOR2HS $T=533820 416760 0 180 $X=528240 $Y=411340
X2231 1374 1408 1399 2 1 XOR2HS $T=537540 457080 0 0 $X=537540 $Y=456700
X2232 1387 1411 1421 2 1 XOR2HS $T=540640 416760 1 0 $X=540640 $Y=411340
X2233 1387 1400 1429 2 1 XOR2HS $T=541880 416760 0 0 $X=541880 $Y=416380
X2234 1457 1436 1442 2 1 XOR2HS $T=554280 426840 1 180 $X=548700 $Y=426460
X2235 1463 1437 1475 2 1 XOR2HS $T=551800 497400 0 0 $X=551800 $Y=497020
X2236 1466 1437 1477 2 1 XOR2HS $T=552420 507480 0 0 $X=552420 $Y=507100
X2237 1457 1406 1455 2 1 XOR2HS $T=559240 426840 0 180 $X=553660 $Y=421420
X2238 1403 1460 1502 2 1 XOR2HS $T=559240 406680 0 0 $X=559240 $Y=406300
X2239 1434 1479 1510 2 1 XOR2HS $T=560480 426840 0 0 $X=560480 $Y=426460
X2240 1466 1401 1523 2 1 XOR2HS $T=562340 507480 1 0 $X=562340 $Y=502060
X2241 1384 1483 1526 2 1 XOR2HS $T=563580 457080 0 0 $X=563580 $Y=456700
X2242 1438 1487 1544 2 1 XOR2HS $T=567920 507480 1 0 $X=567920 $Y=502060
X2243 1519 1400 1554 2 1 XOR2HS $T=571020 416760 0 0 $X=571020 $Y=416380
X2244 1519 1439 1547 2 1 XOR2HS $T=577840 426840 1 180 $X=572260 $Y=426460
X2245 1506 1557 1571 2 1 XOR2HS $T=574120 467160 1 0 $X=574120 $Y=461740
X2246 1461 1408 1581 2 1 XOR2HS $T=575980 487320 1 0 $X=575980 $Y=481900
X2247 1439 1460 1589 2 1 XOR2HS $T=577840 406680 0 0 $X=577840 $Y=406300
X2248 1461 1413 1590 2 1 XOR2HS $T=577840 477240 0 0 $X=577840 $Y=476860
X2249 1457 1400 1593 2 1 XOR2HS $T=578460 426840 1 0 $X=578460 $Y=421420
X2250 1582 1403 1594 2 1 XOR2HS $T=579080 436920 1 0 $X=579080 $Y=431500
X2251 1411 1460 1597 2 1 XOR2HS $T=580320 416760 1 0 $X=580320 $Y=411340
X2252 1556 1408 1599 2 1 XOR2HS $T=580320 527640 1 0 $X=580320 $Y=522220
X2253 1582 1411 1606 2 1 XOR2HS $T=581560 447000 0 0 $X=581560 $Y=446620
X2254 1556 1388 1611 2 1 XOR2HS $T=582800 497400 0 0 $X=582800 $Y=497020
X2255 1582 1400 1610 2 1 XOR2HS $T=583420 447000 1 0 $X=583420 $Y=441580
X2256 1582 134 1609 2 1 XOR2HS $T=583420 457080 1 0 $X=583420 $Y=451660
X2257 1582 1384 1621 2 1 XOR2HS $T=584660 477240 1 0 $X=584660 $Y=471820
X2258 1601 1571 1639 2 1 XOR2HS $T=589000 467160 1 0 $X=589000 $Y=461740
X2259 1614 1416 1645 2 1 XOR2HS $T=590860 467160 0 0 $X=590860 $Y=466780
X2260 1548 1480 1655 2 1 XOR2HS $T=594580 447000 1 0 $X=594580 $Y=441580
X2261 1658 1639 1670 2 1 XOR2HS $T=597680 477240 1 0 $X=597680 $Y=471820
X2262 1661 1588 1658 2 1 XOR2HS $T=598300 467160 0 0 $X=598300 $Y=466780
X2263 1558 1653 1698 2 1 XOR2HS $T=604500 517560 1 0 $X=604500 $Y=512140
X2264 1673 1655 1705 2 1 XOR2HS $T=606360 447000 1 0 $X=606360 $Y=441580
X2265 1570 1699 1709 2 1 XOR2HS $T=606980 426840 0 0 $X=606980 $Y=426460
X2266 1656 1643 1715 2 1 XOR2HS $T=608220 497400 0 0 $X=608220 $Y=497020
X2267 1645 1706 1721 2 1 XOR2HS $T=609460 477240 1 0 $X=609460 $Y=471820
X2268 1671 1684 1736 2 1 XOR2HS $T=613800 527640 1 0 $X=613800 $Y=522220
X2269 1700 1757 1773 2 1 XOR2HS $T=625580 447000 1 0 $X=625580 $Y=441580
X2270 1565 1721 1775 2 1 XOR2HS $T=626200 477240 1 0 $X=626200 $Y=471820
X2271 1732 1790 1804 2 1 XOR2HS $T=634880 517560 0 0 $X=634880 $Y=517180
X2272 1833 1858 1870 2 1 XOR2HS $T=650380 497400 1 0 $X=650380 $Y=491980
X2273 1853 1795 1871 2 1 XOR2HS $T=650380 507480 0 0 $X=650380 $Y=507100
X2274 1867 1848 1880 2 1 XOR2HS $T=652860 487320 1 0 $X=652860 $Y=481900
X2275 1879 1872 1884 2 1 XOR2HS $T=655340 447000 0 0 $X=655340 $Y=446620
X2276 223 1895 1904 2 1 XOR2HS $T=664640 396600 0 0 $X=664640 $Y=396220
X2277 1914 1916 1922 2 1 XOR2HS $T=670220 457080 1 0 $X=670220 $Y=451660
X2278 1886 1899 1939 2 1 XOR2HS $T=675180 436920 1 0 $X=675180 $Y=431500
X2279 1944 246 1934 2 1 XOR2HS $T=681380 406680 1 180 $X=675800 $Y=406300
X2280 1958 1927 1955 2 1 XOR2HS $T=685720 416760 0 180 $X=680140 $Y=411340
X2281 1958 1898 254 2 1 XOR2HS $T=683860 406680 0 0 $X=683860 $Y=406300
X2282 1966 1899 1978 2 1 XOR2HS $T=683860 447000 0 0 $X=683860 $Y=446620
X2283 1973 1952 1986 2 1 XOR2HS $T=685720 487320 0 0 $X=685720 $Y=486940
X2284 1899 1973 1998 2 1 XOR2HS $T=688820 497400 1 0 $X=688820 $Y=491980
X2285 1973 1932 2008 2 1 XOR2HS $T=690060 487320 1 0 $X=690060 $Y=481900
X2286 222 2003 2014 2 1 XOR2HS $T=691920 406680 1 0 $X=691920 $Y=401260
X2287 250 1932 2013 2 1 XOR2HS $T=691920 436920 0 0 $X=691920 $Y=436540
X2288 1932 1972 2017 2 1 XOR2HS $T=691920 467160 1 0 $X=691920 $Y=461740
X2289 2003 224 2046 2 1 XOR2HS $T=696260 396600 0 0 $X=696260 $Y=396220
X2290 1994 1897 2063 2 1 XOR2HS $T=698740 447000 1 0 $X=698740 $Y=441580
X2291 265 1891 2069 2 1 XOR2HS $T=701220 406680 1 0 $X=701220 $Y=401260
X2292 1895 265 2075 2 1 XOR2HS $T=702460 396600 0 0 $X=702460 $Y=396220
X2293 1973 1897 2092 2 1 XOR2HS $T=704940 477240 1 0 $X=704940 $Y=471820
X2294 251 2031 2076 2 1 XOR2HS $T=711140 426840 1 180 $X=705560 $Y=426460
X2295 1973 1915 2102 2 1 XOR2HS $T=706800 467160 1 0 $X=706800 $Y=461740
X2296 271 272 2113 2 1 XOR2HS $T=709280 396600 1 0 $X=709280 $Y=391180
X2297 2093 2011 2103 2 1 XOR2HS $T=714860 487320 1 180 $X=709280 $Y=486940
X2298 273 1895 276 2 1 XOR2HS $T=711140 396600 0 0 $X=711140 $Y=396220
X2299 2111 1891 2144 2 1 XOR2HS $T=713620 426840 1 0 $X=713620 $Y=421420
X2300 2111 251 2147 2 1 XOR2HS $T=714240 436920 0 0 $X=714240 $Y=436540
X2301 2003 1895 2149 2 1 XOR2HS $T=714860 406680 0 0 $X=714860 $Y=406300
X2302 2111 1898 2150 2 1 XOR2HS $T=714860 426840 0 0 $X=714860 $Y=426460
X2303 271 220 2151 2 1 XOR2HS $T=715480 396600 1 0 $X=715480 $Y=391180
X2304 273 1927 2152 2 1 XOR2HS $T=715480 416760 0 0 $X=715480 $Y=416380
X2305 2111 1927 2153 2 1 XOR2HS $T=715480 447000 0 0 $X=715480 $Y=446620
X2306 274 2139 2159 2 1 XOR2HS $T=716720 537720 1 0 $X=716720 $Y=532300
X2307 273 1891 280 2 1 XOR2HS $T=717340 396600 0 0 $X=717340 $Y=396220
X2308 2060 2021 2189 2 1 XOR2HS $T=723540 467160 1 0 $X=723540 $Y=461740
X2309 2176 2194 2204 2 1 XOR2HS $T=726020 497400 0 0 $X=726020 $Y=497020
X2310 2180 2022 2219 2 1 XOR2HS $T=728500 436920 0 0 $X=728500 $Y=436540
X2311 1997 2169 2230 2 1 XOR2HS $T=739660 467160 0 180 $X=734080 $Y=461740
X2312 2230 2216 2249 2 1 XOR2HS $T=734080 477240 1 0 $X=734080 $Y=471820
X2313 2228 2239 289 2 1 XOR2HS $T=734700 527640 0 0 $X=734700 $Y=527260
X2314 2237 2231 2252 2 1 XOR2HS $T=735320 497400 0 0 $X=735320 $Y=497020
X2315 2070 2209 2272 2 1 XOR2HS $T=739040 426840 1 0 $X=739040 $Y=421420
X2316 2197 2263 2295 2 1 XOR2HS $T=743380 447000 1 0 $X=743380 $Y=441580
X2317 2118 2196 2302 2 1 XOR2HS $T=744620 426840 1 0 $X=744620 $Y=421420
X2318 2219 2131 2303 2 1 XOR2HS $T=744620 447000 0 0 $X=744620 $Y=446620
X2319 2218 2297 2311 2 1 XOR2HS $T=745860 527640 1 0 $X=745860 $Y=522220
X2320 2271 2208 2316 2 1 XOR2HS $T=747100 416760 0 0 $X=747100 $Y=416380
X2321 2317 2312 2329 2 1 XOR2HS $T=750200 527640 0 0 $X=750200 $Y=527260
X2322 2319 2327 2340 2 1 XOR2HS $T=752060 487320 1 0 $X=752060 $Y=481900
X2323 2235 2303 2347 2 1 XOR2HS $T=752680 457080 1 0 $X=752680 $Y=451660
X2324 2323 2244 2330 2 1 XOR2HS $T=759500 436920 1 180 $X=753920 $Y=436540
X2325 2355 2348 2374 2 1 XOR2HS $T=759500 527640 0 0 $X=759500 $Y=527260
X2326 2382 2372 2394 2 1 XOR2HS $T=763840 477240 0 0 $X=763840 $Y=476860
X2327 2243 2360 2404 2 1 XOR2HS $T=766940 416760 0 0 $X=766940 $Y=416380
X2328 2385 2425 2447 2 1 XOR2HS $T=775620 517560 0 0 $X=775620 $Y=517180
X2329 2436 2451 2463 2 1 XOR2HS $T=779340 396600 1 0 $X=779340 $Y=391180
X2330 2473 2468 2488 2 1 XOR2HS $T=784300 447000 0 0 $X=784300 $Y=446620
X2331 2485 2461 2492 2 1 XOR2HS $T=786160 527640 1 0 $X=786160 $Y=522220
X2332 2486 2480 2494 2 1 XOR2HS $T=786780 517560 1 0 $X=786780 $Y=512140
X2333 2491 2487 2501 2 1 XOR2HS $T=788640 436920 0 0 $X=788640 $Y=436540
X2334 2460 2475 2509 2 1 XOR2HS $T=790500 507480 0 0 $X=790500 $Y=507100
X2335 2603 2573 2624 2 1 XOR2HS $T=819640 487320 0 0 $X=819640 $Y=486940
X2336 2639 2638 2696 2 1 XOR2HS $T=837000 447000 1 0 $X=837000 $Y=441580
X2337 2739 2742 2753 2 1 XOR2HS $T=854360 527640 0 0 $X=854360 $Y=527260
X2338 2713 2747 2761 2 1 XOR2HS $T=856840 517560 0 0 $X=856840 $Y=517180
X2339 2795 2766 2808 2 1 XOR2HS $T=871720 487320 0 0 $X=871720 $Y=486940
X2340 2845 2864 2874 2 1 XOR2HS $T=886600 517560 0 0 $X=886600 $Y=517180
X2341 2862 2853 2879 2 1 XOR2HS $T=887840 497400 1 0 $X=887840 $Y=491980
X2342 2881 2867 2892 2 1 XOR2HS $T=891560 507480 1 0 $X=891560 $Y=502060
X2343 2921 2927 2954 2 1 XOR2HS $T=907060 507480 1 0 $X=907060 $Y=502060
X2344 2974 2980 2990 2 1 XOR2HS $T=914500 517560 1 0 $X=914500 $Y=512140
X2345 3019 2964 3039 2 1 XOR2HS $T=924420 537720 1 0 $X=924420 $Y=532300
X2346 3030 2988 3044 2 1 XOR2HS $T=926280 527640 1 0 $X=926280 $Y=522220
X2347 3046 2992 3057 2 1 XOR2HS $T=931860 517560 0 0 $X=931860 $Y=517180
X2348 756 776 1 767 788 691 2 MOAI1S $T=374480 487320 0 0 $X=374480 $Y=486940
X2349 815 834 1 825 824 723 2 MOAI1S $T=387500 487320 1 180 $X=383780 $Y=486940
X2350 835 815 1 844 841 830 2 MOAI1S $T=386260 497400 1 0 $X=386260 $Y=491980
X2351 839 867 1 882 844 880 2 MOAI1S $T=394320 517560 0 0 $X=394320 $Y=517180
X2352 967 937 1 918 974 976 2 MOAI1S $T=414160 507480 1 0 $X=414160 $Y=502060
X2353 904 888 1 790 989 990 2 MOAI1S $T=418500 487320 1 0 $X=418500 $Y=481900
X2354 937 1001 1 956 1026 1022 2 MOAI1S $T=429040 447000 1 0 $X=429040 $Y=441580
X2355 937 1043 1 956 975 1063 2 MOAI1S $T=435240 447000 1 0 $X=435240 $Y=441580
X2356 1059 1044 1 989 1053 1078 2 MOAI1S $T=439580 487320 1 0 $X=439580 $Y=481900
X2357 79 1154 1 1083 1150 71 2 MOAI1S $T=461900 396600 0 180 $X=458180 $Y=391180
X2358 1178 1199 1 1225 1221 1234 2 MOAI1S $T=476160 467160 0 0 $X=476160 $Y=466780
X2359 1337 1333 1 1331 1330 1329 2 MOAI1S $T=517700 416760 1 180 $X=513980 $Y=416380
X2360 1373 1378 1 1367 1376 1370 2 MOAI1S $T=532580 426840 1 180 $X=528860 $Y=426460
X2361 1446 1455 1 1449 1462 148 2 MOAI1S $T=549940 416760 1 0 $X=549940 $Y=411340
X2362 1446 1478 1 1462 1459 152 2 MOAI1S $T=557380 416760 0 180 $X=553660 $Y=411340
X2363 1534 1623 1 1627 1595 1642 2 MOAI1S $T=587760 517560 0 0 $X=587760 $Y=517180
X2364 1889 1925 1 234 1909 1919 2 MOAI1S $T=673940 406680 1 0 $X=673940 $Y=401260
X2365 256 2013 1 1981 2004 1999 2 MOAI1S $T=696260 447000 0 180 $X=692540 $Y=441580
X2366 1994 1992 1 1996 2065 2082 2 MOAI1S $T=703700 457080 0 0 $X=703700 $Y=456700
X2367 2138 2102 1 2104 2161 2169 2 MOAI1S $T=717960 457080 0 0 $X=717960 $Y=456700
X2368 399 2873 1 2866 2860 2844 2 MOAI1S $T=890940 527640 0 180 $X=887220 $Y=522220
X2369 2875 397 1 2866 2865 2829 2 MOAI1S $T=890940 527640 1 180 $X=887220 $Y=527260
X2370 2808 2873 1 2866 2855 2843 2 MOAI1S $T=891560 497400 1 180 $X=887840 $Y=497020
X2371 2863 2833 1 2863 2871 2870 2 MOAI1S $T=892800 426840 0 180 $X=889080 $Y=421420
X2372 2849 404 1 2884 2866 2904 2 MOAI1S $T=895280 517560 1 0 $X=895280 $Y=512140
X2373 2863 2903 1 2863 2895 2893 2 MOAI1S $T=899620 426840 0 180 $X=895900 $Y=421420
X2374 2774 404 1 2907 2899 2914 2 MOAI1S $T=897760 487320 0 0 $X=897760 $Y=486940
X2375 2787 404 1 2896 2907 2943 2 MOAI1S $T=901480 497400 1 0 $X=901480 $Y=491980
X2376 404 2954 1 2972 416 2984 2 MOAI1S $T=912020 497400 1 0 $X=912020 $Y=491980
X2377 2958 2971 1 2863 2967 2962 2 MOAI1S $T=916980 426840 0 180 $X=913260 $Y=421420
X2378 2873 2990 1 3054 3055 3047 2 MOAI1S $T=932480 517560 1 0 $X=932480 $Y=512140
X2379 2873 3044 1 3055 3057 3064 2 MOAI1S $T=932480 527640 1 0 $X=932480 $Y=522220
X2380 3133 3083 1 3123 438 2958 2 MOAI1S $T=959140 426840 0 180 $X=955420 $Y=421420
X2381 3154 3112 1 3137 441 3133 2 MOAI1S $T=961620 416760 1 180 $X=957900 $Y=416380
X2382 3210 3175 1 2958 3217 3220 2 MOAI1S $T=984560 426840 0 0 $X=984560 $Y=426460
X2383 3221 3214 1 3223 3226 3154 2 MOAI1S $T=988900 416760 0 0 $X=988900 $Y=416380
X2384 455 3215 1 3222 3229 3221 2 MOAI1S $T=991380 507480 1 0 $X=991380 $Y=502060
X2385 3210 3231 1 3210 3234 3237 2 MOAI1S $T=995100 436920 0 0 $X=995100 $Y=436540
X2386 3210 3249 1 3210 3245 3227 2 MOAI1S $T=1002540 457080 0 180 $X=998820 $Y=451660
X2387 463 3239 1 3253 468 3255 2 MOAI1S $T=1004400 537720 1 0 $X=1004400 $Y=532300
X2388 3253 3236 1 3253 3262 3246 2 MOAI1S $T=1011220 517560 0 180 $X=1007500 $Y=512140
X2389 3253 3265 1 3253 3270 3243 2 MOAI1S $T=1014940 477240 0 180 $X=1011220 $Y=471820
X2390 515 556 512 2 1 ND2S $T=306280 537720 1 0 $X=306280 $Y=532300
X2391 593 33 32 2 1 ND2S $T=346580 537720 1 180 $X=344720 $Y=537340
X2392 627 643 656 2 1 ND2S $T=348440 436920 0 0 $X=348440 $Y=436540
X2393 656 678 645 2 1 ND2S $T=352780 436920 0 0 $X=352780 $Y=436540
X2394 709 717 38 2 1 ND2S $T=362080 537720 0 0 $X=362080 $Y=537340
X2395 745 655 740 2 1 ND2S $T=365800 517560 0 0 $X=365800 $Y=517180
X2396 43 793 752 2 1 ND2S $T=377580 537720 1 180 $X=375720 $Y=537340
X2397 51 985 53 2 1 ND2S $T=415400 537720 1 0 $X=415400 $Y=532300
X2398 996 992 1005 2 1 ND2S $T=424080 467160 0 0 $X=424080 $Y=466780
X2399 1066 1090 1038 2 1 ND2S $T=445780 457080 1 0 $X=445780 $Y=451660
X2400 811 1114 1101 2 1 ND2S $T=449500 477240 0 0 $X=449500 $Y=476860
X2401 68 1124 1055 2 1 ND2S $T=451980 416760 1 0 $X=451980 $Y=411340
X2402 1154 1083 1160 2 1 ND2S $T=459420 396600 0 0 $X=459420 $Y=396220
X2403 1127 1166 1057 2 1 ND2S $T=459420 477240 0 0 $X=459420 $Y=476860
X2404 1078 1188 1186 2 1 ND2S $T=468100 457080 1 180 $X=466240 $Y=456700
X2405 1192 1150 80 2 1 ND2S $T=469340 396600 1 0 $X=469340 $Y=391180
X2406 4 1266 1236 2 1 ND2S $T=486080 497400 1 0 $X=486080 $Y=491980
X2407 1374 1379 1401 2 1 ND2S $T=533820 436920 0 0 $X=533820 $Y=436540
X2408 1640 1647 1598 2 1 ND2S $T=597060 497400 1 180 $X=595200 $Y=497020
X2409 1657 1684 1667 2 1 ND2S $T=603880 527640 0 180 $X=602020 $Y=522220
X2410 1666 1758 1634 2 1 ND2S $T=621240 487320 0 180 $X=619380 $Y=481900
X2411 1816 1867 1806 2 1 ND2S $T=651000 477240 1 180 $X=649140 $Y=476860
X2412 1828 1879 1832 2 1 ND2S $T=656580 447000 1 0 $X=656580 $Y=441580
X2413 1889 229 1897 2 1 ND2S $T=665260 426840 1 0 $X=665260 $Y=421420
X2414 2006 2020 2026 2 1 ND2S $T=695020 497400 0 0 $X=695020 $Y=497020
X2415 2019 2026 2058 2 1 ND2S $T=698120 497400 1 0 $X=698120 $Y=491980
X2416 2227 2239 2205 2 1 ND2S $T=734700 527640 1 0 $X=734700 $Y=522220
X2417 2241 2237 2221 2 1 ND2S $T=737180 487320 1 180 $X=735320 $Y=486940
X2418 2310 2306 2232 2 1 ND2S $T=749580 517560 1 180 $X=747720 $Y=517180
X2419 2335 2355 2259 2 1 ND2S $T=756400 527640 0 0 $X=756400 $Y=527260
X2420 2377 2385 2342 2 1 ND2S $T=764460 517560 1 180 $X=762600 $Y=517180
X2421 2375 2397 2389 2 1 ND2S $T=767560 527640 1 180 $X=765700 $Y=527260
X2422 2368 2410 2414 2 1 ND2S $T=768800 457080 0 0 $X=768800 $Y=456700
X2423 2392 2408 2318 2 1 ND2S $T=770660 517560 1 180 $X=768800 $Y=517180
X2424 2411 2460 2417 2 1 ND2S $T=776240 507480 0 180 $X=774380 $Y=502060
X2425 302 2437 2424 2 1 ND2S $T=776860 406680 0 180 $X=775000 $Y=401260
X2426 2482 2486 2381 2 1 ND2S $T=788020 507480 0 0 $X=788020 $Y=507100
X2427 2556 2552 2518 2 1 ND2S $T=810340 487320 0 180 $X=808480 $Y=481900
X2428 2562 2557 2540 2 1 ND2S $T=811580 477240 0 180 $X=809720 $Y=471820
X2429 2568 2577 2524 2 1 ND2S $T=812820 477240 1 180 $X=810960 $Y=476860
X2430 2584 2583 2549 2 1 ND2S $T=815920 467160 1 180 $X=814060 $Y=466780
X2431 2599 2607 2554 2 1 ND2S $T=819020 447000 0 180 $X=817160 $Y=441580
X2432 2589 2596 2610 2 1 ND2S $T=818400 426840 1 0 $X=818400 $Y=421420
X2433 2633 2639 2586 2 1 ND2S $T=825840 426840 1 180 $X=823980 $Y=426460
X2434 2616 2631 2600 2 1 ND2S $T=827080 467160 0 180 $X=825220 $Y=461740
X2435 2630 2641 2643 2 1 ND2S $T=826460 416760 0 0 $X=826460 $Y=416380
X2436 2616 2645 2605 2 1 ND2S $T=828940 467160 1 180 $X=827080 $Y=466780
X2437 2647 2659 2616 2 1 ND2S $T=830180 467160 0 180 $X=828320 $Y=461740
X2438 2635 2658 2662 2 1 ND2S $T=830180 416760 0 0 $X=830180 $Y=416380
X2439 2661 2664 2587 2 1 ND2S $T=831420 436920 0 0 $X=831420 $Y=436540
X2440 2677 2685 2544 2 1 ND2S $T=837000 457080 1 0 $X=837000 $Y=451660
X2441 2714 2713 2708 2 1 ND2S $T=845060 517560 1 180 $X=843200 $Y=517180
X2442 2715 2739 2703 2 1 ND2S $T=853120 527640 1 180 $X=851260 $Y=527260
X2443 2752 2760 2744 2 1 ND2S $T=858080 487320 0 180 $X=856220 $Y=481900
X2444 2758 2765 2767 2 1 ND2S $T=861180 507480 1 0 $X=861180 $Y=502060
X2445 2767 2776 2778 2 1 ND2S $T=864900 497400 0 0 $X=864900 $Y=497020
X2446 2794 2795 2726 2 1 ND2S $T=870480 487320 1 180 $X=868620 $Y=486940
X2447 2793 2802 2786 2 1 ND2S $T=872340 517560 0 180 $X=870480 $Y=512140
X2448 2824 2826 2834 2 1 ND2S $T=879780 487320 0 0 $X=879780 $Y=486940
X2449 2835 2845 2812 2 1 ND2S $T=882260 517560 1 180 $X=880400 $Y=517180
X2450 2846 2831 381 2 1 ND2S $T=880400 527640 0 0 $X=880400 $Y=527260
X2451 379 2850 2846 2 1 ND2S $T=881020 537720 0 0 $X=881020 $Y=537340
X2452 2856 2860 2753 2 1 ND2S $T=885980 527640 1 180 $X=884120 $Y=527260
X2453 2861 2862 2816 2 1 ND2S $T=887220 497400 0 180 $X=885360 $Y=491980
X2454 2874 2884 2885 2 1 ND2S $T=892180 517560 1 0 $X=892180 $Y=512140
X2455 2882 2881 2807 2 1 ND2S $T=893420 507480 0 0 $X=893420 $Y=507100
X2456 2879 2896 2885 2 1 ND2S $T=894040 497400 1 0 $X=894040 $Y=491980
X2457 2892 2894 2885 2 1 ND2S $T=898380 497400 1 180 $X=896520 $Y=497020
X2458 2942 2957 2883 2 1 ND2S $T=911400 477240 0 180 $X=909540 $Y=471820
X2459 2932 2974 2935 2 1 ND2S $T=914500 517560 0 180 $X=912640 $Y=512140
X2460 2982 2994 2968 2 1 ND2S $T=916980 497400 0 0 $X=916980 $Y=497020
X2461 2926 3017 2910 2 1 ND2S $T=922560 527640 0 180 $X=920700 $Y=522220
X2462 2996 3026 2952 2 1 ND2S $T=923180 467160 1 180 $X=921320 $Y=466780
X2463 2987 3019 2995 2 1 ND2S $T=923800 537720 0 180 $X=921940 $Y=532300
X2464 3001 3030 3017 2 1 ND2S $T=925660 527640 0 180 $X=923800 $Y=522220
X2465 3004 3035 3020 2 1 ND2S $T=926900 467160 1 0 $X=926900 $Y=461740
X2466 3008 3036 3016 2 1 ND2S $T=928760 517560 0 180 $X=926900 $Y=512140
X2467 3042 3046 3027 2 1 ND2S $T=931240 517560 1 180 $X=929380 $Y=517180
X2468 3089 3109 433 2 1 ND2S $T=951700 537720 0 180 $X=949840 $Y=532300
X2469 3136 3141 3065 2 1 ND2S $T=959140 527640 1 180 $X=957280 $Y=527260
X2470 3131 3116 3130 2 1 ND2S $T=957900 487320 1 0 $X=957900 $Y=481900
X2471 3135 3128 3145 2 1 ND2S $T=958520 467160 0 0 $X=958520 $Y=466780
X2472 3147 3142 443 2 1 ND2S $T=960380 507480 0 0 $X=960380 $Y=507100
X2473 3144 3146 3098 2 1 ND2S $T=963480 497400 1 180 $X=961620 $Y=497020
X2474 3159 3139 3148 2 1 ND2S $T=963480 477240 1 0 $X=963480 $Y=471820
X2475 3168 3156 3157 2 1 ND2S $T=965960 507480 0 0 $X=965960 $Y=507100
X2476 3185 3172 3149 2 1 ND2S $T=967200 497400 0 0 $X=967200 $Y=497020
X2477 3201 3183 3191 2 1 ND2S $T=976500 497400 0 0 $X=976500 $Y=497020
X2478 894 870 1 874 869 843 2 MOAI1H $T=399900 447000 1 180 $X=392460 $Y=446620
X2479 927 1013 1 1007 858 927 2 MOAI1H $T=430280 497400 0 180 $X=422840 $Y=491980
X2480 1164 1158 1 1131 1122 1128 2 MOAI1H $T=462520 447000 1 180 $X=455080 $Y=446620
X2481 1373 1358 1 1366 1361 1359 2 MOAI1H $T=531960 406680 1 180 $X=524520 $Y=406300
X2482 1446 1442 1 1460 1383 1462 2 MOAI1H $T=548080 416760 0 0 $X=548080 $Y=416380
X2483 1482 1473 1 1492 1506 1498 2 MOAI1H $T=557380 467160 1 0 $X=557380 $Y=461740
X2484 1537 1547 1 1550 1570 1546 2 MOAI1H $T=571640 436920 1 0 $X=571640 $Y=431500
X2485 1608 1581 1 1541 1634 1498 2 MOAI1H $T=585280 487320 0 0 $X=585280 $Y=486940
X2486 1608 1590 1 1622 1643 1498 2 MOAI1H $T=587140 477240 0 0 $X=587140 $Y=476860
X2487 1608 1598 1 1647 1656 1498 2 MOAI1H $T=592100 497400 1 0 $X=592100 $Y=491980
X2488 1942 1950 1 1957 1968 1950 2 MOAI1H $T=678900 477240 1 0 $X=678900 $Y=471820
X2489 1925 1955 1 1990 1995 2007 2 MOAI1H $T=686340 416760 1 0 $X=686340 $Y=411340
X2490 2038 2017 1 2041 2068 1985 2 MOAI1H $T=698120 467160 1 0 $X=698120 $Y=461740
X2491 281 2163 1 2160 2196 2034 2 MOAI1H $T=722300 426840 0 0 $X=722300 $Y=426460
X2492 2181 2101 1 2197 2260 2268 2 MOAI1H $T=734700 436920 1 0 $X=734700 $Y=431500
X2493 2271 2208 1 2298 2337 2345 2 MOAI1H $T=748960 416760 1 0 $X=748960 $Y=411340
X2494 2360 2243 1 2376 2379 2349 2 MOAI1H $T=759500 416760 0 0 $X=759500 $Y=416380
X2495 570 557 1 2 INV2 $T=326740 487320 1 180 $X=324880 $Y=486940
X2496 567 568 1 2 INV2 $T=327360 487320 1 0 $X=327360 $Y=481900
X2497 582 577 1 2 INV2 $T=336040 497400 1 180 $X=334180 $Y=497020
X2498 635 597 1 2 INV2 $T=344100 447000 1 180 $X=342240 $Y=446620
X2499 824 842 1 2 INV2 $T=386880 487320 0 180 $X=385020 $Y=481900
X2500 842 843 1 2 INV2 $T=387500 487320 1 0 $X=387500 $Y=481900
X2501 858 815 1 2 INV2 $T=391220 467160 1 180 $X=389360 $Y=466780
X2502 851 794 1 2 INV2 $T=391840 436920 1 180 $X=389980 $Y=436540
X2503 842 844 1 2 INV2 $T=391220 497400 1 0 $X=391220 $Y=491980
X2504 848 824 1 2 INV2 $T=422840 477240 0 0 $X=422840 $Y=476860
X2505 790 952 1 2 INV2 $T=424080 487320 0 0 $X=424080 $Y=486940
X2506 995 1018 1 2 INV2 $T=429660 457080 1 0 $X=429660 $Y=451660
X2507 1039 864 1 2 INV2 $T=435240 467160 1 180 $X=433380 $Y=466780
X2508 1041 927 1 2 INV2 $T=435860 487320 0 180 $X=434000 $Y=481900
X2509 1029 1051 1 2 INV2 $T=435240 436920 1 0 $X=435240 $Y=431500
X2510 1006 888 1 2 INV2 $T=437100 507480 0 180 $X=435240 $Y=502060
X2511 1039 1041 1 2 INV2 $T=437100 477240 1 0 $X=437100 $Y=471820
X2512 1060 790 1 2 INV2 $T=439580 477240 0 0 $X=439580 $Y=476860
X2513 1041 1065 1 2 INV2 $T=440200 477240 1 0 $X=440200 $Y=471820
X2514 1073 1039 1 2 INV2 $T=443920 477240 0 180 $X=442060 $Y=471820
X2515 1162 1181 1 2 INV2 $T=463760 447000 1 0 $X=463760 $Y=441580
X2516 81 949 1 2 INV2 $T=466240 436920 1 180 $X=464380 $Y=436540
X2517 1165 1170 1 2 INV2 $T=465000 416760 0 0 $X=465000 $Y=416380
X2518 1353 1374 1 2 INV2 $T=525760 457080 0 0 $X=525760 $Y=456700
X2519 1385 1353 1 2 INV2 $T=532580 457080 1 180 $X=530720 $Y=456700
X2520 1389 1390 1 2 INV2 $T=532580 457080 0 0 $X=532580 $Y=456700
X2521 1381 1389 1 2 INV2 $T=533200 477240 1 0 $X=533200 $Y=471820
X2522 1374 1415 1 2 INV2 $T=540020 436920 0 180 $X=538160 $Y=431500
X2523 1415 1387 1 2 INV2 $T=541260 426840 0 180 $X=539400 $Y=421420
X2524 1415 1378 1 2 INV2 $T=540640 426840 0 0 $X=540640 $Y=426460
X2525 1390 1373 1 2 INV2 $T=541260 436920 1 0 $X=541260 $Y=431500
X2526 143 1308 1 2 INV2 $T=547460 537720 1 180 $X=545600 $Y=537340
X2527 1451 1462 1 2 INV2 $T=554900 436920 0 0 $X=554900 $Y=436540
X2528 1463 1483 1 2 INV2 $T=561100 487320 1 0 $X=561100 $Y=481900
X2529 1503 1446 1 2 INV2 $T=563580 416760 1 180 $X=561720 $Y=416380
X2530 1503 1482 1 2 INV2 $T=562960 447000 0 0 $X=562960 $Y=446620
X2531 1524 1509 1 2 INV2 $T=567920 447000 0 180 $X=566060 $Y=441580
X2532 1529 1543 1 2 INV2 $T=569780 457080 1 0 $X=569780 $Y=451660
X2533 1529 1549 1 2 INV2 $T=571640 497400 1 0 $X=571640 $Y=491980
X2534 1584 1591 1 2 INV2 $T=580940 517560 1 0 $X=580940 $Y=512140
X2535 1582 1583 1 2 INV2 $T=582800 467160 0 0 $X=582800 $Y=466780
X2536 1595 1602 1 2 INV2 $T=584040 517560 1 0 $X=584040 $Y=512140
X2537 1503 1608 1 2 INV2 $T=591480 477240 1 0 $X=591480 $Y=471820
X2538 1623 1572 1 2 INV2 $T=592720 517560 0 0 $X=592720 $Y=517180
X2539 1364 1648 1 2 INV2 $T=596440 396600 0 0 $X=596440 $Y=396220
X2540 1405 1681 1 2 INV2 $T=603260 426840 0 0 $X=603260 $Y=426460
X2541 1443 1690 1 2 INV2 $T=603260 457080 1 0 $X=603260 $Y=451660
X2542 1428 1677 1 2 INV2 $T=606360 447000 1 180 $X=604500 $Y=446620
X2543 1663 1699 1 2 INV2 $T=610080 426840 0 180 $X=608220 $Y=421420
X2544 1430 1717 1 2 INV2 $T=610700 436920 0 0 $X=610700 $Y=436540
X2545 1689 1755 1 2 INV2 $T=621240 426840 1 0 $X=621240 $Y=421420
X2546 1768 1783 1 2 INV2 $T=628680 497400 1 0 $X=628680 $Y=491980
X2547 1729 1788 1 2 INV2 $T=635500 457080 1 0 $X=635500 $Y=451660
X2548 1789 1842 1 2 INV2 $T=639220 507480 1 0 $X=639220 $Y=502060
X2549 1815 1819 1 2 INV2 $T=641080 497400 1 0 $X=641080 $Y=491980
X2550 1795 1852 1 2 INV2 $T=651000 507480 1 0 $X=651000 $Y=502060
X2551 1889 1913 1 2 INV2 $T=672080 436920 0 180 $X=670220 $Y=431500
X2552 1937 1930 1 2 INV2 $T=678280 426840 1 180 $X=676420 $Y=426460
X2553 243 1894 1 2 INV2 $T=678280 537720 0 180 $X=676420 $Y=532300
X2554 1934 237 1 2 INV2 $T=678900 396600 1 180 $X=677040 $Y=396220
X2555 1902 1958 1 2 INV2 $T=680760 416760 0 0 $X=680760 $Y=416380
X2556 1970 255 1 2 INV2 $T=686340 436920 0 0 $X=686340 $Y=436540
X2557 255 1992 1 2 INV2 $T=689440 447000 1 0 $X=689440 $Y=441580
X2558 1950 1972 1 2 INV2 $T=690680 467160 0 0 $X=690680 $Y=466780
X2559 256 1996 1 2 INV2 $T=693780 447000 0 0 $X=693780 $Y=446620
X2560 1968 2028 1 2 INV2 $T=696260 467160 0 0 $X=696260 $Y=466780
X2561 2028 2062 1 2 INV2 $T=699980 436920 0 0 $X=699980 $Y=436540
X2562 2038 267 1 2 INV2 $T=703700 416760 1 180 $X=701840 $Y=416380
X2563 286 2229 1 2 INV2 $T=732840 537720 0 0 $X=732840 $Y=537340
X2564 2249 2279 1 2 INV2 $T=743380 477240 0 0 $X=743380 $Y=476860
X2565 291 2283 1 2 INV2 $T=744620 537720 0 0 $X=744620 $Y=537340
X2566 2291 2274 1 2 INV2 $T=747100 396600 1 180 $X=745240 $Y=396220
X2567 2285 2290 1 2 INV2 $T=745240 487320 1 0 $X=745240 $Y=481900
X2568 2288 2323 1 2 INV2 $T=749580 436920 1 0 $X=749580 $Y=431500
X2569 2106 2345 1 2 INV2 $T=753920 406680 0 0 $X=753920 $Y=406300
X2570 2300 2343 1 2 INV2 $T=755780 467160 0 0 $X=755780 $Y=466780
X2571 2428 2332 1 2 INV2 $T=776240 497400 0 180 $X=774380 $Y=491980
X2572 2479 2428 1 2 INV2 $T=783680 487320 1 180 $X=781820 $Y=486940
X2573 2483 324 1 2 INV2 $T=804140 396600 0 180 $X=802280 $Y=391180
X2574 2483 2469 1 2 INV2 $T=807860 426840 1 0 $X=807860 $Y=421420
X2575 370 2735 1 2 INV2 $T=859320 537720 1 180 $X=857460 $Y=537340
X2576 2745 2858 1 2 INV2 $T=884740 517560 1 0 $X=884740 $Y=512140
X2577 2911 395 1 2 INV2 $T=900860 406680 1 180 $X=899000 $Y=406300
X2578 2922 2911 1 2 INV2 $T=903960 406680 1 180 $X=902100 $Y=406300
X2579 952 898 1 2 BUF2 $T=411060 487320 1 180 $X=407960 $Y=486940
X2580 941 918 1 2 BUF2 $T=411060 497400 0 180 $X=407960 $Y=491980
X2581 45 978 1 2 BUF2 $T=411680 537720 1 0 $X=411680 $Y=532300
X2582 956 941 1 2 BUF2 $T=416020 447000 1 180 $X=412920 $Y=446620
X2583 973 958 1 2 BUF2 $T=422220 477240 1 180 $X=419120 $Y=476860
X2584 995 973 1 2 BUF2 $T=424080 457080 0 180 $X=420980 $Y=451660
X2585 952 1010 1 2 BUF2 $T=425940 487320 0 0 $X=425940 $Y=486940
X2586 1018 975 1 2 BUF2 $T=431520 457080 1 0 $X=431520 $Y=451660
X2587 1082 1194 1 2 BUF2 $T=462520 537720 1 0 $X=462520 $Y=532300
X2588 1194 1253 1 2 BUF2 $T=481740 527640 1 0 $X=481740 $Y=522220
X2589 1253 1282 1 2 BUF2 $T=489800 497400 1 0 $X=489800 $Y=491980
X2590 116 112 1 2 BUF2 $T=518940 527640 0 180 $X=515840 $Y=522220
X2591 1377 1386 1 2 BUF2 $T=533820 497400 0 0 $X=533820 $Y=497020
X2592 1417 1377 1 2 BUF2 $T=544360 517560 1 0 $X=544360 $Y=512140
X2593 1417 116 1 2 BUF2 $T=546840 527640 0 0 $X=546840 $Y=527260
X2594 1456 1460 1 2 BUF2 $T=552420 436920 1 0 $X=552420 $Y=431500
X2595 1462 1497 1 2 BUF2 $T=557380 416760 1 0 $X=557380 $Y=411340
X2596 1525 1417 1 2 BUF2 $T=570400 527640 1 180 $X=567300 $Y=527260
X2597 1556 1466 1 2 BUF2 $T=574740 517560 0 180 $X=571640 $Y=512140
X2598 167 1525 1 2 BUF2 $T=574740 537720 1 0 $X=574740 $Y=532300
X2599 1583 1500 1 2 BUF2 $T=580320 457080 0 0 $X=580320 $Y=456700
X2600 1619 1580 1 2 BUF2 $T=590860 447000 1 0 $X=590860 $Y=441580
X2601 198 195 1 2 BUF2 $T=642940 406680 0 0 $X=642940 $Y=406300
X2602 212 1837 1 2 BUF2 $T=655340 537720 0 180 $X=652240 $Y=532300
X2603 1885 215 1 2 BUF2 $T=660300 416760 0 180 $X=657200 $Y=411340
X2604 1837 206 1 2 BUF2 $T=657200 537720 1 0 $X=657200 $Y=532300
X2605 1886 1889 1 2 BUF2 $T=667740 436920 0 180 $X=664640 $Y=431500
X2606 1890 1896 1 2 BUF2 $T=669600 467160 0 0 $X=669600 $Y=466780
X2607 1896 1885 1 2 BUF2 $T=673940 436920 1 180 $X=670840 $Y=436540
X2608 1894 240 1 2 BUF2 $T=682620 527640 0 180 $X=679520 $Y=522220
X2609 240 1892 1 2 BUF2 $T=680760 517560 1 0 $X=680760 $Y=512140
X2610 1892 1890 1 2 BUF2 $T=682000 507480 1 0 $X=682000 $Y=502060
X2611 237 1974 1 2 BUF2 $T=685100 396600 0 0 $X=685100 $Y=396220
X2612 1950 1940 1 2 BUF2 $T=688200 467160 1 180 $X=685100 $Y=466780
X2613 234 1990 1 2 BUF2 $T=688820 426840 0 0 $X=688820 $Y=426460
X2614 1972 2031 1 2 BUF2 $T=695640 447000 0 0 $X=695640 $Y=446620
X2615 1969 2038 1 2 BUF2 $T=696880 477240 1 0 $X=696880 $Y=471820
X2616 2062 264 1 2 BUF2 $T=702460 396600 0 180 $X=699360 $Y=391180
X2617 267 2044 1 2 BUF2 $T=702460 426840 0 0 $X=702460 $Y=426460
X2618 2029 2107 1 2 BUF2 $T=709280 477240 0 0 $X=709280 $Y=476860
X2619 2133 271 1 2 BUF2 $T=715480 406680 1 0 $X=715480 $Y=401260
X2620 1992 281 1 2 BUF2 $T=720440 436920 0 0 $X=720440 $Y=436540
X2621 2138 2195 1 2 BUF2 $T=728500 436920 1 0 $X=728500 $Y=431500
X2622 2520 2479 1 2 BUF2 $T=799800 507480 0 180 $X=796700 $Y=502060
X2623 322 2520 1 2 BUF2 $T=807860 517560 1 0 $X=807860 $Y=512140
X2624 2560 322 1 2 BUF2 $T=810960 517560 1 180 $X=807860 $Y=517180
X2625 346 2560 1 2 BUF2 $T=829560 527640 1 180 $X=826460 $Y=527260
X2626 358 355 1 2 BUF2 $T=844440 396600 0 180 $X=841340 $Y=391180
X2627 355 372 1 2 BUF2 $T=862420 396600 0 0 $X=862420 $Y=396220
X2628 2785 2797 1 2 BUF2 $T=889700 467160 0 180 $X=886600 $Y=461740
X2629 2900 2890 1 2 BUF2 $T=897140 457080 0 180 $X=894040 $Y=451660
X2630 2907 2866 1 2 BUF2 $T=900240 497400 0 180 $X=897140 $Y=491980
X2631 2890 2950 1 2 BUF2 $T=906440 436920 0 0 $X=906440 $Y=436540
X2632 2953 2900 1 2 BUF2 $T=910160 477240 1 180 $X=907060 $Y=476860
X2633 3003 2922 1 2 BUF2 $T=923180 406680 1 180 $X=920080 $Y=406300
X2634 2950 3034 1 2 BUF2 $T=921940 447000 1 0 $X=921940 $Y=441580
X2635 3034 3003 1 2 BUF2 $T=938680 416760 1 180 $X=935580 $Y=416380
X2636 431 3081 1 2 BUF2 $T=949220 527640 0 0 $X=949220 $Y=527260
X2637 440 434 1 2 BUF2 $T=957900 396600 0 180 $X=954800 $Y=391180
X2638 2953 3171 1 2 BUF2 $T=964720 477240 0 0 $X=964720 $Y=476860
X2639 3173 3163 1 2 BUF2 $T=974640 447000 0 180 $X=971540 $Y=441580
X2640 3163 3161 1 2 BUF2 $T=975260 426840 0 180 $X=972160 $Y=421420
X2641 451 3194 1 2 BUF2 $T=988280 527640 0 0 $X=988280 $Y=527260
X2642 3250 3291 1 2 BUF2 $T=1024860 507480 1 0 $X=1024860 $Y=502060
X2643 3291 3311 1 2 BUF2 $T=1030440 507480 1 0 $X=1030440 $Y=502060
X2644 3311 3297 1 2 BUF2 $T=1033540 507480 1 180 $X=1030440 $Y=507100
X2645 483 480 1 2 BUF2 $T=1039120 487320 0 180 $X=1036020 $Y=481900
X2646 482 476 1 2 BUF2 $T=1039120 537720 0 180 $X=1036020 $Y=532300
X2647 3336 475 1 2 BUF2 $T=1044700 406680 0 180 $X=1041600 $Y=401260
X2648 3297 3335 1 2 BUF2 $T=1043460 517560 1 0 $X=1043460 $Y=512140
X2649 3330 3350 1 2 BUF2 $T=1067640 447000 0 180 $X=1064540 $Y=441580
X2650 3364 3336 1 2 BUF2 $T=1067020 406680 1 0 $X=1067020 $Y=401260
X2651 3350 3393 1 2 BUF2 $T=1070120 447000 1 0 $X=1070120 $Y=441580
X2652 3395 3368 1 2 BUF2 $T=1073840 477240 0 180 $X=1070740 $Y=471820
X2653 3393 3364 1 2 BUF2 $T=1074460 416760 1 180 $X=1071360 $Y=416380
X2654 3335 3386 1 2 BUF2 $T=1083140 517560 1 0 $X=1083140 $Y=512140
X2655 3395 3422 1 2 BUF2 $T=1091820 477240 1 0 $X=1091820 $Y=471820
X2656 3395 3439 1 2 BUF2 $T=1092440 477240 0 0 $X=1092440 $Y=476860
X2657 3446 3428 1 2 BUF2 $T=1109180 457080 0 180 $X=1106080 $Y=451660
X2658 3431 3455 1 2 BUF2 $T=1106700 507480 0 0 $X=1106700 $Y=507100
X2659 496 498 1 2 BUF2 $T=1113520 537720 1 180 $X=1110420 $Y=537340
X2660 3455 3476 1 2 BUF2 $T=1111660 497400 0 0 $X=1111660 $Y=497020
X2661 692 719 712 2 730 739 1 AO22 $T=363320 507480 0 0 $X=363320 $Y=507100
X2662 1457 1456 1 2 INV3 $T=553040 436920 1 180 $X=550560 $Y=436540
X2663 1463 1487 1 2 INV3 $T=558000 497400 0 0 $X=558000 $Y=497020
X2664 1522 1529 1 2 INV3 $T=569160 497400 1 0 $X=569160 $Y=491980
X2665 1907 1929 1 2 INV3 $T=670840 497400 0 0 $X=670840 $Y=497020
X2666 250 246 1 2 INV3 $T=683240 406680 1 0 $X=683240 $Y=401260
X2667 1979 1950 1 2 INV3 $T=687580 487320 1 0 $X=687580 $Y=481900
X2668 2111 2090 1 2 INV3 $T=713000 467160 1 0 $X=713000 $Y=461740
X2669 2483 2510 1 2 INV3 $T=804140 406680 1 0 $X=804140 $Y=401260
X2670 3171 3218 1 2 INV3 $T=985800 467160 0 0 $X=985800 $Y=466780
X2671 3218 3173 1 2 INV3 $T=986420 467160 1 0 $X=986420 $Y=461740
X2672 872 897 1 2 BUF6 $T=396180 457080 1 0 $X=396180 $Y=451660
X2673 1375 1367 1 2 BUF6 $T=530720 447000 0 180 $X=523280 $Y=441580
X2674 1598 1461 1 2 BUF6 $T=585280 487320 1 180 $X=577840 $Y=486940
X2675 3291 3290 1 2 BUF6 $T=1029200 487320 0 0 $X=1029200 $Y=486940
X2676 3393 3419 1 2 BUF6 $T=1098020 426840 0 0 $X=1098020 $Y=426460
X2677 750 1 753 757 669 767 2 OAI22S $T=369520 477240 1 0 $X=369520 $Y=471820
X2678 788 1 753 767 716 750 2 OAI22S $T=377580 477240 1 180 $X=373860 $Y=476860
X2679 801 1 753 766 808 829 2 OAI22S $T=382540 457080 0 0 $X=382540 $Y=456700
X2680 933 1 921 918 845 912 2 OAI22S $T=406720 517560 0 180 $X=403000 $Y=512140
X2681 935 1 953 941 759 943 2 OAI22S $T=412920 457080 0 180 $X=409200 $Y=451660
X2682 963 1 953 951 736 941 2 OAI22S $T=412920 467160 1 180 $X=409200 $Y=466780
X2683 960 1 921 957 961 941 2 OAI22S $T=416020 497400 0 180 $X=412300 $Y=491980
X2684 974 1 921 918 965 962 2 OAI22S $T=417880 517560 1 180 $X=414160 $Y=517180
X2685 886 1 753 925 991 1020 2 OAI22S $T=422840 457080 0 0 $X=422840 $Y=456700
X2686 1040 1 925 753 1031 1020 2 OAI22S $T=435860 457080 1 180 $X=432140 $Y=456700
X2687 1113 1 1104 1061 1129 1118 2 OAI22S $T=457560 477240 0 180 $X=453840 $Y=471820
X2688 1376 1 1391 1367 1362 1393 2 OAI22S $T=531960 436920 1 0 $X=531960 $Y=431500
X2689 1402 1 1391 1395 128 1367 2 OAI22S $T=537540 406680 0 180 $X=533820 $Y=401260
X2690 1393 1 1391 1367 1404 1402 2 OAI22S $T=533820 426840 1 0 $X=533820 $Y=421420
X2691 1391 1 1448 1366 1458 1440 2 OAI22S $T=548700 406680 1 0 $X=548700 $Y=401260
X2692 1470 1 1471 1476 1480 1462 2 OAI22S $T=553660 447000 1 0 $X=553660 $Y=441580
X2693 1524 1 1530 1543 1531 1507 2 OAI22S $T=570400 467160 1 0 $X=570400 $Y=461740
X2694 1546 1 1524 1552 1548 1543 2 OAI22S $T=575980 447000 0 180 $X=572260 $Y=441580
X2695 1542 1 1535 1550 1553 1567 2 OAI22S $T=572880 406680 0 0 $X=572880 $Y=406300
X2696 1524 1 1544 1549 1558 1562 2 OAI22S $T=572880 507480 0 0 $X=572880 $Y=507100
X2697 1909 1 237 234 235 230 2 OAI22S $T=673320 396600 0 180 $X=669600 $Y=391180
X2698 1974 1 2040 1990 2033 1913 2 OAI22S $T=700600 436920 0 180 $X=696880 $Y=431500
X2699 2044 1 2051 2041 2061 2052 2 OAI22S $T=699360 457080 1 0 $X=699360 $Y=451660
X2700 1985 1 2044 2041 2056 2023 2 OAI22S $T=704320 477240 0 180 $X=700600 $Y=471820
X2701 2083 1 2044 2062 2067 2051 2 OAI22S $T=706800 436920 1 180 $X=703080 $Y=436540
X2702 270 1 267 264 2081 2084 2 OAI22S $T=704320 396600 1 0 $X=704320 $Y=391180
X2703 508 2 5 7 507 1 9 FA1S $T=287060 537720 0 0 $X=287060 $Y=537340
X2704 1332 2 1346 1328 1362 1 1337 FA1S $T=511500 436920 1 0 $X=511500 $Y=431500
X2705 2064 2 2085 2053 2012 1 2110 FA1S $T=698120 517560 0 0 $X=698120 $Y=517180
X2706 2143 2 2105 1964 2098 1 2200 FA1S $T=712380 517560 0 0 $X=712380 $Y=517180
X2707 2183 2 2172 2032 2112 1 2224 FA1S $T=720440 517560 1 0 $X=720440 $Y=512140
X2708 2255 2 2233 2024 2234 1 2296 FA1S $T=734700 517560 1 0 $X=734700 $Y=512140
X2709 2328 2 2320 1963 2309 1 2341 FA1S $T=748960 507480 0 0 $X=748960 $Y=507100
X2710 2339 2 2315 1956 2367 1 2373 FA1S $T=750820 507480 1 0 $X=750820 $Y=502060
X2711 2396 2 2351 1910 2420 1 2393 FA1S $T=763220 487320 0 0 $X=763220 $Y=486940
X2712 2474 2 2452 1901 2484 1 2498 FA1S $T=780580 477240 0 0 $X=780580 $Y=476860
X2713 2478 2 2489 2453 2493 1 2502 FA1S $T=781200 487320 1 0 $X=781200 $Y=481900
X2714 2490 2 2457 2466 2462 1 2511 FA1S $T=784300 467160 0 0 $X=784300 $Y=466780
X2715 2526 2 321 2537 2519 1 2500 FA1S $T=805380 447000 0 180 $X=793600 $Y=441580
X2716 2527 2 2515 2541 2531 1 2506 FA1S $T=805380 457080 0 180 $X=793600 $Y=451660
X2717 2528 2 2513 2533 2514 1 2503 FA1S $T=805380 457080 1 180 $X=793600 $Y=456700
X2718 2529 2 2538 1905 2532 1 2504 FA1S $T=805380 467160 0 180 $X=793600 $Y=461740
X2719 2525 2 320 319 2508 1 2547 FA1S $T=796080 426840 1 0 $X=796080 $Y=421420
X2720 2543 2 2559 1893 2548 1 2578 FA1S $T=801040 426840 0 0 $X=801040 $Y=426460
X2721 2558 2 333 326 2569 1 2604 FA1S $T=806000 416760 1 0 $X=806000 $Y=411340
X2722 2563 2 330 2516 2555 1 2572 FA1S $T=807240 416760 0 0 $X=807240 $Y=416380
X2723 2580 2 332 2523 2553 1 2618 FA1S $T=809720 406680 1 0 $X=809720 $Y=401260
X2724 2594 2 336 335 2581 1 2614 FA1S $T=813440 406680 0 0 $X=813440 $Y=406300
X2725 2673 2 2682 349 350 1 351 FA1S $T=829560 537720 1 0 $X=829560 $Y=532300
X2726 2707 2 2687 356 2689 1 2720 FA1S $T=838240 497400 1 0 $X=838240 $Y=491980
X2727 2728 2 2681 362 2705 1 2741 FA1S $T=845060 507480 1 0 $X=845060 $Y=502060
X2728 2748 2 2730 365 2634 1 2755 FA1S $T=851880 527640 1 0 $X=851880 $Y=522220
X2729 2764 2 2722 368 2593 1 2779 FA1S $T=856220 537720 1 0 $X=856220 $Y=532300
X2730 2872 2 2871 2833 2827 1 3491 FA1S $T=885360 416760 0 0 $X=885360 $Y=416380
X2731 2901 2 2837 409 2653 1 2926 FA1S $T=892800 517560 0 0 $X=892800 $Y=517180
X2732 2910 2 2828 406 2671 1 2937 FA1S $T=895900 537720 0 0 $X=895900 $Y=537340
X2733 2915 2 2823 411 1941 1 2938 FA1S $T=896520 507480 0 0 $X=896520 $Y=507100
X2734 2919 2 2895 2903 2872 1 3492 FA1S $T=897760 416760 0 0 $X=897760 $Y=416380
X2735 2977 2 2967 2971 2919 1 3493 FA1S $T=911400 416760 0 0 $X=911400 $Y=416380
X2736 3213 2 3217 3175 2977 1 3494 FA1S $T=980840 436920 1 0 $X=980840 $Y=431500
X2737 3242 2 3234 3231 3213 1 3495 FA1S $T=994480 436920 1 0 $X=994480 $Y=431500
X2738 3248 2 3262 3236 3242 1 3496 FA1S $T=1006880 517560 1 180 $X=995100 $Y=517180
X2739 3251 2 468 3239 3248 1 3497 FA1S $T=1006880 527640 0 180 $X=995100 $Y=522220
X2740 467 2 3270 3265 3261 1 3498 FA1S $T=1011220 477240 0 180 $X=999440 $Y=471820
X2741 3261 2 3245 3249 3251 1 3499 FA1S $T=1005020 477240 0 0 $X=1005020 $Y=476860
X2742 890 882 1 2 INV4 $T=399900 507480 1 180 $X=396800 $Y=507100
X2743 882 872 1 2 INV4 $T=398660 497400 0 0 $X=398660 $Y=497020
X2744 1170 1236 1 2 INV4 $T=477400 487320 0 0 $X=477400 $Y=486940
X2745 1236 1369 1 2 INV4 $T=527620 517560 0 180 $X=524520 $Y=512140
X2746 1929 1973 1 2 INV4 $T=685100 497400 1 0 $X=685100 $Y=491980
X2747 3275 3267 1 2 INV4 $T=1024240 436920 0 180 $X=1021140 $Y=431500
X2748 3298 3238 1 2 INV4 $T=1026720 447000 1 0 $X=1026720 $Y=441580
X2749 3290 3378 1 2 INV4 $T=1054000 487320 0 0 $X=1054000 $Y=486940
X2750 3378 3402 1 2 INV4 $T=1084380 487320 0 0 $X=1084380 $Y=486940
X2751 1184 1192 80 79 1 2 NR3HP $T=469960 396600 1 180 $X=462520 $Y=396220
X2752 1065 1066 1 1054 2 OR2T $T=439580 457080 1 0 $X=439580 $Y=451660
X2753 1003 1155 1 1197 2 OR2T $T=461900 436920 1 0 $X=461900 $Y=431500
X2754 2249 2226 1 2236 2 OR2T $T=740280 477240 1 180 $X=734080 $Y=476860
X2755 2254 2245 1 2286 2 OR2T $T=740280 457080 0 0 $X=740280 $Y=456700
X2756 865 1028 1012 1027 2 864 1 AOI13HS $T=431520 477240 0 0 $X=431520 $Y=476860
X2757 1356 1469 1433 1472 2 1463 1 AOI13HS $T=553040 477240 0 0 $X=553040 $Y=476860
X2758 1953 2 1928 246 1954 1 NR3 $T=683860 447000 1 180 $X=680760 $Y=446620
X2759 1065 1061 1086 1 2 1110 OA12 $T=448260 487320 1 0 $X=448260 $Y=481900
X2760 1085 1061 1114 1 2 1152 OA12 $T=452600 477240 0 0 $X=452600 $Y=476860
X2761 1130 1123 1149 1 2 1168 OA12 $T=459420 507480 0 0 $X=459420 $Y=507100
X2762 1255 1240 1248 1 2 1262 OA12 $T=482360 487320 0 0 $X=482360 $Y=486940
X2763 1397 1375 1410 1 2 1416 OA12 $T=535060 467160 1 0 $X=535060 $Y=461740
X2764 1549 1487 1561 1 2 1568 OA12 $T=574120 497400 1 0 $X=574120 $Y=491980
X2765 1795 1776 1789 1 2 1807 OA12 $T=636740 507480 0 0 $X=636740 $Y=507100
X2766 1991 1990 2009 1 2 2022 OA12 $T=691920 436920 1 0 $X=691920 $Y=431500
X2767 1950 1968 2037 1 2 2048 OA12 $T=696260 487320 1 0 $X=696260 $Y=481900
X2768 2000 2035 2026 1 2 2049 OA12 $T=696880 497400 0 0 $X=696880 $Y=497020
X2769 2108 274 275 1 2 2136 OA12 $T=712380 537720 1 0 $X=712380 $Y=532300
X2770 2231 2247 2221 1 2 2278 OA12 $T=739660 497400 1 0 $X=739660 $Y=491980
X2771 2664 2638 2656 1 2 2695 OA12 $T=835760 436920 0 0 $X=835760 $Y=436540
X2772 2916 2782 2905 1 2 2887 OA12 $T=901480 537720 0 180 $X=897760 $Y=532300
X2773 3011 419 2999 1 2 2907 OA12 $T=921940 497400 0 180 $X=918220 $Y=491980
X2774 3093 3094 3095 1 2 422 OA12 $T=947980 477240 0 0 $X=947980 $Y=476860
X2775 3093 3094 3095 1 2 2931 OA12 $T=947980 487320 1 0 $X=947980 $Y=481900
X2776 3088 3113 3090 1 2 3095 OA12 $T=952940 477240 1 0 $X=952940 $Y=471820
X2777 3093 3094 3095 1 2 436 OA12 $T=952940 477240 0 0 $X=952940 $Y=476860
X2778 3093 3094 3095 1 2 414 OA12 $T=952940 487320 1 0 $X=952940 $Y=481900
X2779 921 912 1 918 859 905 2 OAI22H $T=407960 507480 1 180 $X=400520 $Y=507100
X2780 1359 1390 1 1367 1405 1412 2 OAI22H $T=531340 447000 1 0 $X=531340 $Y=441580
X2781 1391 1412 1 1409 1430 1418 2 OAI22H $T=538780 447000 1 0 $X=538780 $Y=441580
X2782 1418 1390 1 1409 1428 1419 2 OAI22H $T=538780 447000 0 0 $X=538780 $Y=446620
X2783 1535 1510 1 1550 168 1542 2 OAI22H $T=569780 416760 1 0 $X=569780 $Y=411340
X2784 1975 1974 1 242 2001 1989 2 OAI22H $T=688200 396600 0 0 $X=688200 $Y=396220
X2785 2007 1974 1 1990 2039 2047 2 OAI22H $T=693780 416760 1 0 $X=693780 $Y=411340
X2786 563 8 24 28 1 2 QDFFRBP $T=324260 537720 1 0 $X=324260 $Y=532300
X2787 704 8 608 36 1 2 QDFFRBP $T=372620 527640 1 180 $X=360220 $Y=527260
X2788 49 8 45 890 1 2 QDFFRBP $T=409820 537720 0 180 $X=397420 $Y=532300
X2789 988 8 949 995 1 2 QDFFRBP $T=420980 416760 0 0 $X=420980 $Y=416380
X2790 1034 61 978 1073 1 2 QDFFRBP $T=433380 517560 1 0 $X=433380 $Y=512140
X2791 1037 61 1050 1060 1 2 QDFFRBP $T=434000 426840 1 0 $X=434000 $Y=421420
X2792 1241 66 1212 922 1 2 QDFFRBP $T=481120 517560 1 180 $X=468720 $Y=517180
X2793 1687 159 173 1516 1 2 QDFFRBP $T=603880 537720 0 180 $X=591480 $Y=532300
X2794 180 159 173 1598 1 2 QDFFRBP $T=605120 537720 1 180 $X=592720 $Y=537340
X2795 1881 204 1890 1907 1 2 QDFFRBP $T=657200 497400 0 0 $X=657200 $Y=497020
X2796 218 204 1896 1908 1 2 QDFFRBP $T=657820 457080 1 0 $X=657820 $Y=451660
X2797 1883 204 1888 1928 1 2 QDFFRBP $T=657820 477240 1 0 $X=657820 $Y=471820
X2798 238 204 1885 1886 1 2 QDFFRBP $T=673940 447000 0 180 $X=661540 $Y=441580
X2799 231 204 1888 1916 1 2 QDFFRBP $T=667740 477240 0 0 $X=667740 $Y=476860
X2800 2463 204 318 2515 1 2 QDFFRBP $T=788020 396600 0 0 $X=788020 $Y=396220
X2801 1850 204 2510 2541 1 2 QDFFRBP $T=794840 416760 0 0 $X=794840 $Y=416380
X2802 1310 61 1287 2 1 920 QDFFRBS $T=507160 517560 0 180 $X=495380 $Y=512140
X2803 1452 66 1467 2 1 1388 QDFFRBS $T=549320 517560 0 0 $X=549320 $Y=517180
X2804 160 159 1525 2 1 1563 QDFFRBS $T=562960 527640 1 0 $X=562960 $Y=522220
X2805 1294 1308 1 1300 1313 2 101 1249 105 OAI222S $T=504060 537720 1 0 $X=504060 $Y=532300
X2806 99 1308 1 102 1313 2 94 1238 105 OAI222S $T=509640 537720 1 0 $X=509640 $Y=532300
X2807 118 1308 1 107 1313 2 119 1241 105 OAI222S $T=520180 527640 0 0 $X=520180 $Y=527260
X2808 125 1308 1 1314 1313 2 1360 1310 105 OAI222S $T=529480 527640 0 180 $X=523900 $Y=522220
X2809 145 101 1 1294 149 2 150 1452 153 OAI222S $T=549320 537720 0 0 $X=549320 $Y=537340
X2810 145 1360 1 125 149 2 156 1488 153 OAI222S $T=563580 537720 1 180 $X=558000 $Y=537340
X2811 1367 2 1 1366 BUF3 $T=530100 406680 0 180 $X=526380 $Y=401260
X2812 1461 2 1 1356 BUF3 $T=555520 487320 0 180 $X=551800 $Y=481900
X2813 1462 2 1 1498 BUF3 $T=559240 447000 0 0 $X=559240 $Y=446620
X2814 3161 2 1 3204 BUF3 $T=978360 406680 0 0 $X=978360 $Y=406300
X2815 3431 2 1 3395 BUF3 $T=1094920 487320 0 180 $X=1091200 $Y=481900
X2816 3467 2 1 3446 BUF3 $T=1125920 447000 0 0 $X=1125920 $Y=446620
X2817 1369 117 1 2 INV6 $T=527620 517560 1 0 $X=527620 $Y=512140
X2818 3204 3271 1 2 INV6 $T=1014320 406680 1 180 $X=1009360 $Y=406300
X2819 3271 3276 1 2 INV6 $T=1014940 406680 0 0 $X=1014940 $Y=406300
X2820 3276 3275 1 2 INV6 $T=1015560 416760 0 0 $X=1015560 $Y=416380
X2821 3267 3298 1 2 INV6 $T=1025480 447000 0 180 $X=1020520 $Y=441580
X2822 3454 3467 1 2 INV6 $T=1106080 436920 1 0 $X=1106080 $Y=431500
X2823 857 1 865 2 BUF4CK $T=392460 497400 0 0 $X=392460 $Y=497020
X2824 127 1 1313 2 BUF4CK $T=531340 537720 1 180 $X=526380 $Y=537340
X2825 1461 1 1457 2 BUF4CK $T=554280 447000 1 180 $X=549320 $Y=446620
X2826 1516 1 1463 2 BUF4CK $T=572880 487320 0 0 $X=572880 $Y=486940
X2827 1913 1 1900 2 BUF4CK $T=672080 426840 1 180 $X=667120 $Y=426460
X2828 1908 1 250 2 BUF4CK $T=680760 436920 1 0 $X=680760 $Y=431500
X2829 1973 1 2111 2 BUF4CK $T=708660 467160 0 0 $X=708660 $Y=466780
X2830 243 1 2483 2 BUF4CK $T=791120 416760 0 180 $X=786160 $Y=411340
X2831 2510 318 1 2 BUF4 $T=803520 396600 0 0 $X=803520 $Y=396220
X2832 3402 3431 1 2 BUF4 $T=1093680 507480 0 180 $X=1089340 $Y=502060
X2833 243 2953 1 2 INV4CK $T=931240 487320 1 0 $X=931240 $Y=481900
X2834 737 723 691 2 1 651 XOR3 $T=367660 487320 1 180 $X=356500 $Y=486940
X2835 851 826 800 2 1 805 XOR3 $T=392460 436920 0 180 $X=381300 $Y=431500
X2836 1153 1179 1129 2 1 1223 XOR3 $T=465000 487320 0 0 $X=465000 $Y=486940
X2837 522 517 526 519 1 2 ND3P $T=312480 497400 1 180 $X=307520 $Y=497020
X2838 537 525 538 531 1 2 ND3P $T=318060 487320 1 180 $X=313100 $Y=486940
X2839 552 522 530 543 1 2 ND3P $T=323020 497400 1 180 $X=318060 $Y=497020
X2840 555 548 559 550 1 2 ND3P $T=324260 517560 0 180 $X=319300 $Y=512140
X2841 552 537 564 541 1 2 ND3P $T=326120 487320 0 180 $X=321160 $Y=481900
X2842 544 555 558 543 1 2 ND3P $T=327360 507480 0 180 $X=322400 $Y=502060
X2843 552 581 543 577 1 2 ND3P $T=325500 497400 0 0 $X=325500 $Y=497020
X2844 581 571 591 576 1 2 ND3P $T=332940 507480 0 180 $X=327980 $Y=502060
X2845 552 594 598 543 1 2 ND3P $T=339140 507480 0 180 $X=334180 $Y=502060
X2846 594 615 605 601 1 2 ND3P $T=334800 517560 1 0 $X=334800 $Y=512140
X2847 1260 1254 1244 1235 1 2 ND3P $T=487940 477240 1 180 $X=482980 $Y=476860
X2848 2218 2256 2283 2253 1 2 ND3P $T=744620 537720 0 180 $X=739660 $Y=532300
X2849 562 607 582 1 2 OR2P $T=340380 497400 1 180 $X=336660 $Y=497020
X2850 1670 1742 1816 1 2 OR2P $T=635500 477240 0 0 $X=635500 $Y=476860
X2851 2199 2211 2241 1 2 OR2P $T=734080 487320 1 0 $X=734080 $Y=481900
X2852 2300 2264 2325 1 2 OR2P $T=749580 477240 1 0 $X=749580 $Y=471820
X2853 2347 2353 2354 1 2 OR2P $T=761980 457080 1 180 $X=758260 $Y=456700
X2854 1798 2 1 1793 1830 NR2F $T=642940 436920 1 180 $X=636120 $Y=436540
X2855 1803 2 1 1797 1834 NR2F $T=639220 416760 0 0 $X=639220 $Y=416380
X2856 1830 2 1 1834 1836 NR2F $T=643560 436920 1 0 $X=643560 $Y=431500
X2857 1747 204 1885 3500 1893 1 2 DFFRBP $T=651620 416760 0 0 $X=651620 $Y=416380
X2858 311 204 2510 2523 3501 1 2 DFFRBP $T=788020 406680 1 0 $X=788020 $Y=401260
X2859 327 232 2479 2508 3502 1 2 DFFRBP $T=806000 497400 0 180 $X=791740 $Y=491980
X2860 323 232 2520 3503 2548 1 2 DFFRBP $T=800420 507480 1 0 $X=800420 $Y=502060
X2861 334 232 2520 2569 3504 1 2 DFFRBP $T=809720 507480 0 0 $X=809720 $Y=507100
X2862 345 232 2520 2581 3505 1 2 DFFRBP $T=826460 517560 0 180 $X=812200 $Y=512140
X2863 925 1 2 806 INV3CK $T=406100 457080 1 180 $X=403000 $Y=456700
X2864 557 546 1 542 534 2 OAI12HP $T=324880 497400 0 180 $X=314340 $Y=491980
X2865 1210 1205 1 1229 1240 2 OAI12HP $T=469340 497400 0 0 $X=469340 $Y=497020
X2866 1471 1498 1 1504 1528 2 OAI12HP $T=557380 457080 1 0 $X=557380 $Y=451660
X2867 1765 1732 1 1756 1795 2 OAI12HP $T=626200 507480 0 0 $X=626200 $Y=507100
X2868 1846 1841 1 1809 1817 2 OAI12HP $T=652240 457080 0 180 $X=641700 $Y=451660
X2869 1928 1940 1 1945 256 2 OAI12HP $T=678900 457080 1 0 $X=678900 $Y=451660
X2870 1507 1524 1 1490 1517 1508 2 OAI112HS $T=569160 487320 0 180 $X=564820 $Y=481900
X2871 514 8 509 10 1 2 3506 DFFRBN $T=311860 517560 0 180 $X=298840 $Y=512140
X2872 524 8 509 11 1 2 3507 DFFRBN $T=311860 517560 1 180 $X=298840 $Y=517180
X2873 521 8 509 14 1 2 3508 DFFRBN $T=316820 527640 0 180 $X=303800 $Y=522220
X2874 758 8 45 46 1 2 3509 DFFRBN $T=377580 537720 1 0 $X=377580 $Y=532300
X2875 1215 66 82 78 1 2 3510 DFFRBN $T=474300 537720 1 180 $X=461280 $Y=537340
X2876 1882 204 1885 1905 1 2 3511 DFFRBN $T=657200 436920 0 0 $X=657200 $Y=436540
X2877 316 232 322 2531 1 2 3512 DFFRBN $T=792980 517560 1 0 $X=792980 $Y=512140
X2878 317 232 322 2519 1 2 3513 DFFRBN $T=792980 517560 0 0 $X=792980 $Y=517180
X2879 342 232 2576 2553 1 2 3514 DFFRBN $T=821500 497400 1 180 $X=808480 $Y=497020
X2880 597 1 604 614 2 544 ND3HT $T=334180 447000 0 0 $X=334180 $Y=446620
X2881 597 1 604 614 2 552 ND3HT $T=334180 457080 1 0 $X=334180 $Y=451660
X2882 613 1 619 633 2 614 ND3HT $T=338520 436920 1 0 $X=338520 $Y=431500
X2883 1163 1 1227 1232 2 633 ND3HT $T=472440 436920 1 0 $X=472440 $Y=431500
X2884 1197 1 1193 1228 2 1232 ND3HT $T=483600 447000 0 180 $X=476160 $Y=441580
X2885 1806 1 1827 1820 2 1835 ND3HT $T=648520 477240 0 180 $X=641080 $Y=471820
X2886 1816 1 1784 1833 2 1820 ND3HT $T=642320 487320 1 0 $X=642320 $Y=481900
X2887 1819 1 1838 1844 2 1833 ND3HT $T=642940 497400 1 0 $X=642940 $Y=491980
X2888 1823 1 1839 1849 2 198 ND3HT $T=643560 426840 1 0 $X=643560 $Y=421420
X2889 1857 1 1836 1835 2 1849 ND3HT $T=651620 447000 0 180 $X=644180 $Y=441580
X2890 2241 1 2236 2258 2 2269 ND3HT $T=745240 487320 0 180 $X=737800 $Y=481900
X2891 292 1 2314 2256 2 2338 ND3HT $T=758260 537720 0 180 $X=750820 $Y=532300
X2892 2325 1 2354 2319 2 2366 ND3HT $T=765080 477240 0 180 $X=757640 $Y=471820
X2893 2384 1 2371 2366 2 2400 ND3HT $T=771280 467160 0 180 $X=763840 $Y=461740
X2894 2430 1 2427 2400 2 2433 ND3HT $T=779960 447000 0 180 $X=772520 $Y=441580
X2895 2426 1 2440 2433 2 304 ND3HT $T=774380 436920 1 0 $X=774380 $Y=431500
X2896 307 1 2448 2338 2 306 ND3HT $T=783680 537720 1 180 $X=776240 $Y=537340
X2897 889 888 702 884 1 885 2 AOI22S $T=399900 477240 0 180 $X=396180 $Y=471820
X2898 904 888 726 887 1 885 2 AOI22S $T=399900 487320 0 180 $X=396180 $Y=481900
X2899 884 888 772 911 1 885 2 AOI22S $T=397420 467160 0 0 $X=397420 $Y=466780
X2900 887 888 725 889 1 885 2 AOI22S $T=399900 477240 1 0 $X=399900 $Y=471820
X2901 911 917 855 913 1 885 2 AOI22S $T=403000 467160 0 0 $X=403000 $Y=466780
X2902 913 917 908 924 1 885 2 AOI22S $T=403620 477240 1 0 $X=403620 $Y=471820
X2903 924 917 914 964 1 944 2 AOI22S $T=412300 477240 1 0 $X=412300 $Y=471820
X2904 964 917 997 1004 1 944 2 AOI22S $T=424080 477240 1 0 $X=424080 $Y=471820
X2905 1044 1059 1081 1069 1 944 2 AOI22S $T=443920 487320 1 180 $X=440200 $Y=486940
X2906 1093 1059 1088 1023 1 65 2 AOI22S $T=448260 497400 0 0 $X=448260 $Y=497020
X2907 65 1116 1146 1059 1 1115 2 AOI22S $T=458800 497400 0 180 $X=455080 $Y=491980
X2908 1512 1580 1586 1536 1 1574 2 AOI22S $T=581560 426840 1 180 $X=577840 $Y=426460
X2909 1594 1580 1604 1610 1 1574 2 AOI22S $T=584660 436920 1 0 $X=584660 $Y=431500
X2910 1521 1574 1632 1536 1 1580 2 AOI22S $T=589000 426840 1 180 $X=585280 $Y=426460
X2911 1477 1602 1612 1534 1 1623 2 AOI22S $T=585900 517560 1 0 $X=585900 $Y=512140
X2912 1609 1619 1614 1621 1 1605 2 AOI22S $T=587140 457080 0 0 $X=587140 $Y=456700
X2913 1577 1619 1624 1606 1 1605 2 AOI22S $T=588380 447000 0 0 $X=588380 $Y=446620
X2914 1606 1619 1629 1609 1 1605 2 AOI22S $T=589000 457080 1 0 $X=589000 $Y=451660
X2915 1611 1619 1631 1523 1 1623 2 AOI22S $T=589000 497400 0 0 $X=589000 $Y=497020
X2916 1521 1580 1638 1594 1 1574 2 AOI22S $T=591480 426840 0 0 $X=591480 $Y=426460
X2917 1998 2054 2050 2057 1 2029 2 AOI22S $T=700600 487320 0 0 $X=700600 $Y=486940
X2918 2008 2054 2093 1986 1 2029 2 AOI22S $T=708660 487320 1 180 $X=704940 $Y=486940
X2919 2102 2054 2134 2092 1 2107 2 AOI22S $T=715480 477240 0 180 $X=711760 $Y=471820
X2920 2147 2153 2175 2138 1 2107 2 AOI22S $T=723540 447000 0 0 $X=723540 $Y=446620
X2921 2147 2107 2180 2150 1 2138 2 AOI22S $T=724160 436920 1 0 $X=724160 $Y=431500
X2922 2046 2195 2207 2113 1 2174 2 AOI22S $T=731600 396600 1 180 $X=727880 $Y=396220
X2923 2144 2195 2210 2150 1 2174 2 AOI22S $T=729740 426840 0 0 $X=729740 $Y=426460
X2924 1023 1 2 1127 BUF1CK $T=452600 487320 1 0 $X=452600 $Y=481900
X2925 1282 1 2 1287 BUF1CK $T=500340 507480 0 180 $X=497860 $Y=502060
X2926 1282 1 2 1286 BUF1CK $T=502200 487320 0 0 $X=502200 $Y=486940
X2927 1282 1 2 1335 BUF1CK $T=515220 487320 1 0 $X=515220 $Y=481900
X2928 1538 1 2 1640 BUF1CK $T=585280 497400 1 0 $X=585280 $Y=491980
X2929 2125 1 2 2138 BUF1CK $T=713620 457080 0 0 $X=713620 $Y=456700
X2930 2856 1 2 2885 BUF1CK $T=891560 527640 1 0 $X=891560 $Y=522220
X2931 699 731 1 742 627 2 OAI12H $T=375100 426840 1 180 $X=368900 $Y=426460
X2932 1353 1357 1 1363 1375 2 OAI12H $T=522660 467160 1 0 $X=522660 $Y=461740
X2933 1396 1366 1 1423 1427 2 OAI12H $T=536920 396600 0 0 $X=536920 $Y=396220
X2934 1526 1543 1 1559 1592 2 OAI12H $T=575980 457080 1 0 $X=575980 $Y=451660
X2935 1728 1733 1 1737 1757 2 OAI12H $T=615040 447000 1 0 $X=615040 $Y=441580
X2936 1750 1778 1 1770 1793 2 OAI12H $T=629300 436920 0 0 $X=629300 $Y=436540
X2937 1781 1755 1 1764 1803 2 OAI12H $T=631160 426840 1 0 $X=631160 $Y=421420
X2938 2052 2044 1 1962 2021 2 OAI12H $T=701840 457080 1 180 $X=695640 $Y=456700
X2939 2121 2034 1 2179 2208 2 OAI12H $T=721680 416760 0 0 $X=721680 $Y=416380
X2940 2176 2201 1 2167 2231 2 OAI12H $T=729120 487320 0 0 $X=729120 $Y=486940
X2941 2222 2223 1 2215 2254 2 OAI12H $T=733460 457080 0 0 $X=733460 $Y=456700
X2942 2368 2380 1 2383 2416 2 OAI12H $T=762600 447000 0 0 $X=762600 $Y=446620
X2943 2375 2398 1 2403 2418 2 OAI12H $T=767560 537720 1 0 $X=767560 $Y=532300
X2944 2693 2700 1 2708 2718 2 OAI12H $T=839480 517560 1 0 $X=839480 $Y=512140
X2945 2821 2745 1 2839 392 2 OAI12H $T=878540 517560 1 0 $X=878540 $Y=512140
X2946 80 1 79 1154 1209 2 ND3S $T=465000 396600 1 0 $X=465000 $Y=391180
X2947 1832 1 1855 1866 1857 2 ND3S $T=655340 447000 0 180 $X=652860 $Y=441580
X2948 1972 1 2042 2037 2038 2 ND3S $T=698120 477240 0 0 $X=698120 $Y=476860
X2949 543 544 2 535 534 1 AOI12H $T=321780 507480 0 180 $X=315580 $Y=502060
X2950 564 544 2 539 549 1 AOI12H $T=326740 477240 1 180 $X=320540 $Y=476860
X2951 586 544 2 569 573 1 AOI12H $T=332940 457080 1 180 $X=326740 $Y=456700
X2952 1707 1722 2 1732 1695 1 AOI12H $T=620000 517560 1 180 $X=613800 $Y=517180
X2953 2126 2049 2 2176 2099 1 AOI12H $T=718580 497400 1 0 $X=718580 $Y=491980
X2954 2424 305 2 2451 2439 1 AOI12H $T=779340 396600 0 0 $X=779340 $Y=396220
X2955 2100 2086 2116 1 2 2127 HA1 $T=706800 527640 1 0 $X=706800 $Y=522220
X2956 2673 2720 2698 1 2 2691 HA1 $T=847540 497400 1 180 $X=839480 $Y=497020
X2957 360 359 2686 1 2 2701 HA1 $T=849400 537720 0 180 $X=841340 $Y=532300
X2958 2748 2779 2800 1 2 2803 HA1 $T=866140 527640 1 0 $X=866140 $Y=522220
X2959 2728 2755 2801 1 2 2798 HA1 $T=868620 507480 0 0 $X=868620 $Y=507100
X2960 2707 2741 2805 1 2 2814 HA1 $T=869860 497400 1 0 $X=869860 $Y=491980
X2961 2764 382 387 1 2 2815 HA1 $T=873580 537720 1 0 $X=873580 $Y=532300
X2962 2920 2915 2944 1 2 2956 HA1 $T=902100 497400 0 0 $X=902100 $Y=497020
X2963 2901 2938 2960 1 2 2993 HA1 $T=910160 507480 0 0 $X=910160 $Y=507100
X2964 2910 2926 3005 1 2 3018 HA1 $T=915120 517560 0 0 $X=915120 $Y=517180
X2965 415 2937 3032 1 2 426 HA1 $T=923800 537720 0 0 $X=923800 $Y=537340
X2966 1048 1 1054 925 2 ND2T $T=434620 457080 1 0 $X=434620 $Y=451660
X2967 283 1 285 2218 2 ND2T $T=727260 537720 0 0 $X=727260 $Y=537340
X2968 2290 1 2269 2319 2 ND2T $T=747100 487320 1 0 $X=747100 $Y=481900
X2969 1822 1812 1850 1845 1 2 MXL2H $T=642320 406680 1 0 $X=642320 $Y=401260
X2970 1930 1900 234 1906 1 2 MXL2H $T=677040 426840 0 180 $X=668360 $Y=421420
X2971 1605 1610 2 1580 1628 1577 1 AOI22H $T=584660 436920 0 0 $X=584660 $Y=436540
X2972 2174 2014 2 2195 284 2046 1 AOI22H $T=723540 406680 1 0 $X=723540 $Y=401260
X2973 2174 2113 2 2151 2213 2195 1 AOI22H $T=725400 406680 0 0 $X=725400 $Y=406300
X2974 2174 2149 2 2195 2209 2144 1 AOI22H $T=725400 426840 1 0 $X=725400 $Y=421420
X2975 2174 2151 2 2195 2220 2149 1 AOI22H $T=727260 416760 1 0 $X=727260 $Y=411340
X2976 1464 1483 1503 1445 1 2 MXL2HP $T=554900 467160 0 0 $X=554900 $Y=466780
X2977 897 936 955 1 2 XNR2H $T=419740 436920 0 180 $X=411060 $Y=431500
X2978 927 848 1014 1 2 XNR2H $T=420360 497400 0 0 $X=420360 $Y=497020
X2979 1352 1391 1356 1 2 XNR2H $T=529480 477240 0 0 $X=529480 $Y=476860
X2980 1444 1451 1487 1 2 XNR2H $T=549940 497400 1 0 $X=549940 $Y=491980
X2981 1630 1653 1659 1 2 XNR2H $T=590860 507480 0 0 $X=590860 $Y=507100
X2982 1649 1666 1675 1 2 XNR2H $T=593960 487320 0 0 $X=593960 $Y=486940
X2983 181 1710 179 1 2 XNR2H $T=604500 396600 1 0 $X=604500 $Y=391180
X2984 1734 1729 1724 1 2 XNR2H $T=622480 457080 1 180 $X=613800 $Y=456700
X2985 1709 1746 1720 1 2 XNR2H $T=615660 426840 0 0 $X=615660 $Y=426460
X2986 1689 1767 1678 1 2 XNR2H $T=621240 436920 1 0 $X=621240 $Y=431500
X2987 1666 1768 1726 1 2 XNR2H $T=634880 487320 1 180 $X=626200 $Y=486940
X2988 1751 1797 1686 1 2 XNR2H $T=643560 416760 0 180 $X=634880 $Y=411340
X2989 2404 2429 2349 1 2 XNR2H $T=783060 416760 1 180 $X=774380 $Y=416380
X2990 607 519 623 576 1 2 OA12P $T=344100 507480 0 180 $X=339760 $Y=502060
X2991 1828 1834 1805 1839 1 2 OA12P $T=643560 426840 0 0 $X=643560 $Y=426460
X2992 2477 2458 2476 2426 1 2 OA12P $T=788020 436920 0 180 $X=783680 $Y=431500
X2993 511 8 509 6 1 2 3515 DFFRBS $T=302560 527640 1 180 $X=289540 $Y=527260
X2994 620 8 608 3516 1 2 26 DFFRBS $T=347200 527640 0 180 $X=334180 $Y=522220
X2995 2148 232 2122 2 1 2105 2097 232 2122 2145 506 ICV_20 $T=710520 507480 1 0 $X=710520 $Y=502060
X2996 2159 232 2122 2 1 2234 2204 232 2122 2172 506 ICV_20 $T=735320 507480 0 180 $X=723540 $Y=502060
X2997 2732 344 2717 2 1 2702 2702 344 2717 2743 506 ICV_20 $T=841960 436920 1 0 $X=841960 $Y=431500
X2998 2888 2813 2890 2 1 2917 2934 2813 2890 2833 506 ICV_20 $T=905200 447000 0 180 $X=893420 $Y=441580
X2999 3070 2813 3063 2 1 3101 3101 2813 3063 3069 506 ICV_20 $T=952320 426840 0 180 $X=940540 $Y=421420
X3000 445 430 3169 2 1 3190 3190 430 3169 3157 506 ICV_20 $T=974640 537720 0 180 $X=962860 $Y=532300
X3001 3247 3151 3250 2 1 3272 3266 3151 3250 3229 506 ICV_20 $T=1010600 507480 0 180 $X=998820 $Y=502060
X3002 3320 3151 3335 2 1 3339 3339 3327 3311 3319 506 ICV_20 $T=1047800 507480 0 180 $X=1036020 $Y=502060
X3003 3326 3327 3311 2 1 3347 3347 3327 3311 3324 506 ICV_20 $T=1050900 497400 0 180 $X=1039120 $Y=491980
X3004 3367 3327 3350 2 1 3342 3343 3327 3350 3367 506 ICV_20 $T=1047800 447000 1 0 $X=1047800 $Y=441580
X3005 3349 3327 3368 2 1 3375 3344 3327 3290 3349 506 ICV_20 $T=1062060 477240 0 180 $X=1050280 $Y=471820
X3006 3360 3327 3330 2 1 3381 3381 485 3330 3361 506 ICV_20 $T=1067640 436920 0 180 $X=1055860 $Y=431500
X3007 3372 485 3336 2 1 3394 488 485 3336 3369 506 ICV_20 $T=1072600 396600 0 180 $X=1060820 $Y=391180
X3008 3452 486 3455 2 1 3472 3477 486 3455 3452 506 ICV_20 $T=1114760 517560 0 180 $X=1102980 $Y=512140
X3009 3462 3327 3446 2 1 3480 3480 3327 3446 3444 506 ICV_20 $T=1123440 447000 0 180 $X=1111660 $Y=441580
X3010 3468 3327 3439 2 1 3481 3481 3327 3428 3463 506 ICV_20 $T=1124060 467160 0 180 $X=1112280 $Y=461740
X3011 3464 3327 3476 2 1 3483 3483 3327 3439 3468 506 ICV_20 $T=1124680 477240 0 180 $X=1112900 $Y=471820
X3012 2870 2857 2 2844 1 396 MUX2S $T=890940 426840 1 180 $X=886600 $Y=426460
X3013 2893 2857 2 2843 1 401 MUX2S $T=897140 426840 1 180 $X=892800 $Y=426460
X3014 2962 2857 2 2914 1 421 MUX2S $T=913260 426840 0 0 $X=913260 $Y=426460
X3015 3220 2857 2 2943 1 458 MUX2S $T=990760 426840 0 0 $X=990760 $Y=426460
X3016 3227 2857 2 449 1 461 MUX2S $T=992000 447000 0 0 $X=992000 $Y=446620
X3017 3243 462 2 447 1 459 MUX2S $T=999440 477240 0 180 $X=995100 $Y=471820
X3018 3255 462 2 445 1 456 MUX2S $T=1000060 537720 1 180 $X=995720 $Y=537340
X3019 3237 462 2 2891 1 465 MUX2S $T=998200 447000 1 0 $X=998200 $Y=441580
X3020 3246 462 2 2904 1 464 MUX2S $T=999440 517560 1 0 $X=999440 $Y=512140
X3021 1143 1192 2 1 1250 1132 MUX2 $T=474920 406680 1 0 $X=474920 $Y=401260
X3022 2841 2857 2 1 384 2829 MUX2 $T=885360 426840 1 180 $X=881020 $Y=426460
X3023 2851 2863 2 1 2841 389 MUX2 $T=887220 426840 0 180 $X=882880 $Y=421420
X3024 2902 2931 2 1 2888 2897 MUX2 $T=902100 467160 0 180 $X=897760 $Y=461740
X3025 2963 422 2 1 2973 2883 MUX2 $T=918220 477240 1 180 $X=913880 $Y=476860
X3026 2978 414 2 1 2998 2952 MUX2 $T=915740 467160 0 0 $X=915740 $Y=466780
X3027 2997 2931 2 1 3022 3020 MUX2 $T=920700 467160 1 0 $X=920700 $Y=461740
X3028 3087 422 2 1 432 433 MUX2 $T=946740 537720 1 180 $X=942400 $Y=537340
X3029 3080 414 2 1 3091 3073 MUX2 $T=944880 467160 1 0 $X=944880 $Y=461740
X3030 3084 436 2 1 3082 3049 MUX2 $T=951700 457080 1 180 $X=947360 $Y=456700
X3031 3110 2931 2 1 3125 3098 MUX2 $T=952940 497400 0 0 $X=952940 $Y=497020
X3032 3138 436 2 1 3114 3086 MUX2 $T=958520 457080 1 180 $X=954180 $Y=456700
X3033 3150 414 2 1 3158 3065 MUX2 $T=967200 527640 1 180 $X=962860 $Y=527260
X3034 3162 436 2 1 3181 3145 MUX2 $T=964720 457080 1 0 $X=964720 $Y=451660
X3035 3165 422 2 1 3178 3148 MUX2 $T=965340 477240 1 0 $X=965340 $Y=471820
X3036 3187 414 2 1 3174 3157 MUX2 $T=973400 527640 1 180 $X=969060 $Y=527260
X3037 3189 436 2 1 3202 3149 MUX2 $T=973400 487320 1 0 $X=973400 $Y=481900
X3038 3193 2931 2 1 3200 3191 MUX2 $T=975260 497400 1 0 $X=975260 $Y=491980
X3039 2727 2735 2 2745 2718 1 AOI12HP $T=859940 517560 0 180 $X=849400 $Y=512140
X3040 1673 1480 1548 1689 1 2 MAO222P $T=600160 447000 1 0 $X=600160 $Y=441580
X3041 1106 1105 1112 2 1 1131 AN3 $T=450120 447000 0 0 $X=450120 $Y=446620
X3042 114 1308 1 110 1313 105 1275 123 2 OAI222H $T=515220 537720 0 0 $X=515220 $Y=537340
X3043 94 1308 1 1313 99 105 1365 126 2 OAI222H $T=517700 537720 1 0 $X=517700 $Y=532300
X3044 1767 1798 1746 1 2 XNR2HP $T=625580 426840 0 0 $X=625580 $Y=426460
X3045 1929 1960 1 2 INV2CK $T=682000 497400 1 0 $X=682000 $Y=491980
X3046 397 2856 1 2 INV2CK $T=890940 527640 0 0 $X=890940 $Y=527260
X3047 95 61 1286 2 1 821 1279 61 1286 1303 506 ICV_22 $T=503440 477240 1 180 $X=491660 $Y=476860
X3048 2699 344 2712 2 1 2732 2734 344 2712 2699 506 ICV_22 $T=840720 447000 0 0 $X=840720 $Y=446620
X3049 2736 344 355 2 1 357 2709 344 355 2736 506 ICV_22 $T=854360 396600 1 180 $X=842580 $Y=396220
X3050 2780 344 355 2 1 2746 2749 344 2770 2780 506 ICV_22 $T=867380 406680 1 180 $X=855600 $Y=406300
X3051 2792 344 372 2 1 2836 2822 344 2770 2792 506 ICV_22 $T=869240 396600 0 0 $X=869240 $Y=396220
X3052 413 391 2922 2 1 2989 2989 391 2922 2930 506 ICV_22 $T=907680 396600 0 0 $X=907680 $Y=396220
X3053 3086 2813 3079 2 1 3102 3102 2813 3079 3138 506 ICV_22 $T=962860 447000 1 180 $X=951080 $Y=446620
X3054 3170 391 3075 2 1 3124 3112 2813 3161 3170 506 ICV_22 $T=968440 406680 1 180 $X=956660 $Y=406300
X3055 3280 3151 3267 2 1 3257 3258 3151 3267 3280 506 ICV_22 $T=1018660 436920 1 180 $X=1006880 $Y=436540
X3056 3285 430 472 2 1 3263 3263 430 472 3287 506 ICV_22 $T=1019900 527640 1 180 $X=1008120 $Y=527260
X3057 3284 3151 3294 2 1 3302 3301 3151 3290 3284 506 ICV_22 $T=1018040 477240 0 0 $X=1018040 $Y=476860
X3058 3288 3151 3238 2 1 3307 3303 3151 3238 3288 506 ICV_22 $T=1019900 447000 0 0 $X=1019900 $Y=446620
X3059 3333 3151 3315 2 1 3354 3354 485 3315 3331 506 ICV_22 $T=1042840 416760 0 0 $X=1042840 $Y=416380
X3060 3340 446 3336 2 1 3372 3365 485 3336 3340 506 ICV_22 $T=1047180 396600 0 0 $X=1047180 $Y=396220
X3061 3382 485 3364 2 1 3362 3361 485 3364 3382 506 ICV_22 $T=1068260 416760 1 180 $X=1056480 $Y=416380
X3062 3413 3327 3368 2 1 3345 3391 3327 3368 3412 506 ICV_22 $T=1081280 457080 1 180 $X=1069500 $Y=456700
X3063 3416 3327 3401 2 1 3435 3434 3327 3401 3416 506 ICV_22 $T=1083140 436920 0 0 $X=1083140 $Y=436540
X3064 3418 485 3419 2 1 3420 3435 3327 3401 3418 506 ICV_22 $T=1083760 426840 0 0 $X=1083760 $Y=426460
X3065 3436 485 3440 2 1 3453 3448 485 3440 3408 506 ICV_22 $T=1094300 396600 0 0 $X=1094300 $Y=396220
X3066 3457 3327 3446 2 1 3441 3444 3327 3428 3457 506 ICV_22 $T=1109180 436920 1 180 $X=1097400 $Y=436540
X3067 3458 3327 3428 2 1 3442 3442 3327 3428 3459 506 ICV_22 $T=1109180 457080 1 180 $X=1097400 $Y=456700
X3068 3473 485 3440 2 1 3448 3451 485 3440 3470 506 ICV_22 $T=1113520 406680 1 180 $X=1101740 $Y=406300
X3069 3449 486 3396 2 1 3450 3450 486 498 3456 506 ICV_22 $T=1113520 527640 1 180 $X=1101740 $Y=527260
X3070 3475 485 3467 2 1 3489 3484 3327 3467 3474 506 ICV_22 $T=1114140 426840 0 0 $X=1114140 $Y=426460
X3071 3478 486 3455 2 1 3486 3487 486 498 3478 506 ICV_22 $T=1116620 517560 0 0 $X=1116620 $Y=517180
X3072 3479 486 498 2 1 3487 3488 486 498 3479 506 ICV_22 $T=1116620 527640 0 0 $X=1116620 $Y=527260
X3073 977 8 949 2 1 931 931 8 949 955 506 ICV_23 $T=419120 416760 0 180 $X=406720 $Y=411340
X3074 1045 61 978 2 1 56 58 8 978 1014 506 ICV_23 $T=434620 527640 0 180 $X=422220 $Y=522220
X3075 1035 61 949 2 1 1080 1094 61 1050 1037 506 ICV_23 $T=433380 416760 1 0 $X=433380 $Y=411340
X3076 124 61 1377 2 1 1411 1407 61 1377 1352 506 ICV_23 $T=525760 507480 1 0 $X=525760 $Y=502060
X3077 2252 232 2122 2 1 2233 2190 232 2122 2309 506 ICV_23 $T=748340 507480 0 180 $X=735940 $Y=502060
X3078 3023 391 2922 2 1 3058 3024 2813 3003 3023 506 ICV_23 $T=924420 406680 1 0 $X=924420 $Y=401260
X3079 3072 391 434 2 1 435 3077 391 429 3072 506 ICV_23 $T=940540 396600 1 0 $X=940540 $Y=391180
X3080 3105 2813 3075 2 1 3074 3069 2813 3063 3105 506 ICV_23 $T=953560 416760 0 180 $X=941160 $Y=411340
X3081 3199 446 3161 2 1 3182 3177 446 3161 3199 506 ICV_23 $T=982080 416760 0 180 $X=969680 $Y=411340
X3082 460 446 450 2 1 3212 3212 446 450 3240 506 ICV_23 $T=996960 396600 0 180 $X=984560 $Y=391180
X3083 466 446 3204 2 1 3226 3233 446 3204 3259 506 ICV_23 $T=1007500 406680 0 180 $X=995100 $Y=401260
X3084 3296 430 476 2 1 3293 3293 430 472 478 506 ICV_23 $T=1033540 537720 0 180 $X=1021140 $Y=532300
X3085 3321 3151 3290 2 1 3344 3346 3327 3290 3321 506 ICV_23 $T=1036640 477240 1 0 $X=1036640 $Y=471820
X3086 3342 3327 3350 2 1 3341 3341 3327 481 3383 506 ICV_23 $T=1059580 457080 0 180 $X=1047180 $Y=451660
X3087 3410 3327 3393 2 1 3388 3388 3327 3401 3411 506 ICV_23 $T=1081280 436920 0 180 $X=1068880 $Y=431500
X3088 3408 485 3417 2 1 3430 3430 485 3417 3407 506 ICV_23 $T=1080040 406680 1 0 $X=1080040 $Y=401260
X3089 3345 3327 3428 2 1 3414 3437 3327 3422 3413 506 ICV_23 $T=1082520 457080 1 0 $X=1082520 $Y=451660
X3090 3412 3327 3422 2 1 3415 3415 3327 3422 3437 506 ICV_23 $T=1094920 467160 0 180 $X=1082520 $Y=461740
X3091 3443 3327 3439 2 1 3460 3460 3327 3439 3445 506 ICV_23 $T=1098020 477240 1 0 $X=1098020 $Y=471820
X3092 135 131 1 1382 2 OR2B1S $T=538160 396600 0 180 $X=535060 $Y=391180
X3093 1971 1925 1 2009 2 OR2B1S $T=691920 426840 0 0 $X=691920 $Y=426460
X3094 2851 389 1 2827 2 OR2B1S $T=883500 416760 1 180 $X=880400 $Y=416380
X3095 310 204 318 2516 1 2 3517 DFFRBT $T=786160 396600 1 0 $X=786160 $Y=391180
X3096 325 204 2469 2559 1 2 2574 DFFRBT $T=802900 436920 1 0 $X=802900 $Y=431500
X3097 1745 159 182 1 2 1556 QDFFRBT $T=620000 537720 0 180 $X=606360 $Y=532300
X3098 308 204 2510 1 2 2537 QDFFRBT $T=789260 406680 0 0 $X=789260 $Y=406300
X3099 2003 2114 1 2 INV1CK $T=714240 406680 1 180 $X=712380 $Y=406300
X3100 1908 1914 1 2 BUF2CK $T=675800 457080 1 0 $X=675800 $Y=451660
X3101 1544 1549 1537 1475 2 1 1518 MAOI1HP $T=575360 497400 1 180 $X=562340 $Y=497020
X3102 1419 1390 1 1409 1443 1441 2 OAI22HP $T=538160 457080 1 0 $X=538160 $Y=451660
X3103 975 980 1 1000 956 975 2 MOAI1HP $T=416640 436920 0 0 $X=416640 $Y=436540
.ENDS
***************************************
.SUBCKT TIE1 O VCC GND
** N=4 EP=3 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OA12S B2 B1 A1 VCC GND O
** N=7 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_25 1 2 3 4 5 7 8 9 10 11 12 14 15 16 17 18 19 20 21 22
+ 24 25 26 27 28 29 30 32 33 34 35 36 37 38 39 40 41 42 43 44
+ 45 46 47 48 49 50 51 52 53 54 56 57 58 59 60 61 62 63 64 65
+ 67 68 69 70 71 72 73 74 75 76 77 78 79 80 82 83 84 85 86 87
+ 88 89 90 91 92 93 94 95 96 97 98 99 100 101 102 103 104 105 106 107
+ 108 109 110 111 112 113 114 115 116 117 118 119 120 121 122 123 124 125 126 127
+ 128 129 130 131 132 133 134 135 136 137 138 139 140 141 142 143 144 146 147 148
+ 149 150 151 152 153 154 155 156 157 158 159 160 161 162 163 164 165 166 167 168
+ 169 170 171 172 173 174 175 176 177 205
** N=1012 EP=170 IP=5185 FDC=0
X0 3 1 2 4 BUF1S $T=231880 225240 0 180 $X=229400 $Y=219820
X1 5 1 2 3 BUF1S $T=334180 225240 0 180 $X=331700 $Y=219820
X2 136 1 2 110 BUF1S $T=887220 225240 0 180 $X=884740 $Y=219820
X3 150 1 2 136 BUF1S $T=929380 225240 0 180 $X=926900 $Y=219820
X4 175 1 2 177 BUF1S $T=1125920 336120 1 0 $X=1125920 $Y=330700
X5 335 2 1 82 BUF1 $T=686340 376440 0 0 $X=686340 $Y=376060
X6 110 2 1 5 BUF1 $T=773140 225240 0 180 $X=770660 $Y=219820
X7 118 2 1 495 BUF1 $T=801040 376440 0 180 $X=798560 $Y=371020
X8 496 2 1 509 BUF1 $T=806000 305880 0 0 $X=806000 $Y=305500
X9 512 2 1 513 BUF1 $T=815300 376440 1 180 $X=812820 $Y=376060
X10 532 2 1 511 BUF1 $T=823980 356280 0 180 $X=821500 $Y=350860
X11 531 2 1 528 BUF1 $T=824600 285720 1 180 $X=822120 $Y=285340
X12 530 2 1 126 BUF1 $T=827700 376440 1 180 $X=825220 $Y=376060
X13 529 2 1 531 BUF1 $T=827700 305880 1 0 $X=827700 $Y=300460
X14 529 2 1 550 BUF1 $T=832040 315960 0 0 $X=832040 $Y=315580
X15 550 2 1 563 BUF1 $T=854360 315960 0 0 $X=854360 $Y=315580
X16 550 2 1 578 BUF1 $T=859320 305880 1 180 $X=856840 $Y=305500
X17 550 2 1 589 BUF1 $T=860560 315960 0 0 $X=860560 $Y=315580
X18 642 2 1 644 BUF1 $T=903960 376440 1 0 $X=903960 $Y=371020
X19 626 2 1 651 BUF1 $T=907060 315960 0 0 $X=907060 $Y=315580
X20 626 2 1 642 BUF1 $T=909540 376440 1 0 $X=909540 $Y=371020
X21 641 2 1 683 BUF1 $T=912020 295800 0 0 $X=912020 $Y=295420
X22 667 2 1 685 BUF1 $T=913260 265560 0 0 $X=913260 $Y=265180
X23 642 2 1 684 BUF1 $T=913880 376440 1 0 $X=913880 $Y=371020
X24 682 2 1 667 BUF1 $T=916980 275640 1 180 $X=914500 $Y=275260
X25 683 2 1 699 BUF1 $T=931860 295800 0 0 $X=931860 $Y=295420
X26 684 2 1 148 BUF1 $T=936200 376440 0 0 $X=936200 $Y=376060
X27 683 2 1 719 BUF1 $T=937440 295800 0 0 $X=937440 $Y=295420
X28 682 2 1 720 BUF1 $T=946740 275640 1 0 $X=946740 $Y=270220
X29 719 2 1 745 BUF1 $T=950460 315960 1 0 $X=950460 $Y=310540
X30 720 2 1 749 BUF1 $T=951080 275640 1 0 $X=951080 $Y=270220
X31 151 2 1 774 BUF1 $T=963480 376440 1 0 $X=963480 $Y=371020
X32 769 2 1 789 BUF1 $T=968440 295800 0 0 $X=968440 $Y=295420
X33 770 2 1 763 BUF1 $T=968440 356280 1 0 $X=968440 $Y=350860
X34 772 2 1 771 BUF1 $T=974640 326040 0 0 $X=974640 $Y=325660
X35 778 2 1 773 BUF1 $T=982080 275640 0 0 $X=982080 $Y=275260
X36 774 2 1 160 BUF1 $T=982080 386520 0 0 $X=982080 $Y=386140
X37 772 2 1 805 BUF1 $T=995720 346200 1 0 $X=995720 $Y=340780
X38 160 2 1 819 BUF1 $T=999440 386520 1 180 $X=996960 $Y=386140
X39 160 2 1 839 BUF1 $T=1001300 386520 0 0 $X=1001300 $Y=386140
X40 830 2 1 824 BUF1 $T=1003160 326040 0 0 $X=1003160 $Y=325660
X41 828 2 1 850 BUF1 $T=1005020 285720 0 0 $X=1005020 $Y=285340
X42 850 2 1 823 BUF1 $T=1008740 275640 1 180 $X=1006260 $Y=275260
X43 823 2 1 856 BUF1 $T=1007500 275640 1 0 $X=1007500 $Y=270220
X44 167 2 1 168 BUF1 $T=1016180 225240 1 0 $X=1016180 $Y=219820
X45 857 2 1 896 BUF1 $T=1027340 356280 1 0 $X=1027340 $Y=350860
X46 853 2 1 901 BUF1 $T=1033540 315960 1 0 $X=1033540 $Y=310540
X47 895 2 1 870 BUF1 $T=1040980 285720 0 0 $X=1040980 $Y=285340
X48 919 2 1 900 BUF1 $T=1044700 346200 0 0 $X=1044700 $Y=345820
X49 919 2 1 922 BUF1 $T=1057720 336120 1 180 $X=1055240 $Y=335740
X50 951 2 1 946 BUF1 $T=1070120 376440 1 0 $X=1070120 $Y=371020
X51 951 2 1 975 BUF1 $T=1080040 366360 0 0 $X=1080040 $Y=365980
X52 974 2 1 994 BUF1 $T=1100500 326040 0 0 $X=1100500 $Y=325660
X53 975 2 1 995 BUF1 $T=1103600 366360 0 0 $X=1103600 $Y=365980
X54 995 2 1 989 BUF1 $T=1106700 376440 0 0 $X=1106700 $Y=376060
X55 176 2 1 150 BUF1 $T=1119720 225240 0 180 $X=1117240 $Y=219820
X56 177 2 1 176 BUF1 $T=1129020 285720 1 180 $X=1126540 $Y=285340
X57 7 8 9 2 1 10 QDFFRBN $T=454460 386520 0 0 $X=454460 $Y=386140
X58 12 8 9 2 1 11 QDFFRBN $T=481120 386520 1 180 $X=469340 $Y=386140
X59 56 58 59 2 1 61 QDFFRBN $T=648520 386520 0 0 $X=648520 $Y=386140
X60 492 58 114 2 1 493 QDFFRBN $T=783060 315960 0 0 $X=783060 $Y=315580
X61 498 58 114 2 1 491 QDFFRBN $T=795460 326040 0 180 $X=783680 $Y=320620
X62 493 58 496 2 1 500 QDFFRBN $T=785540 305880 0 0 $X=785540 $Y=305500
X63 494 58 496 2 1 498 QDFFRBN $T=785540 315960 1 0 $X=785540 $Y=310540
X64 500 502 509 2 1 520 QDFFRBN $T=799800 305880 1 0 $X=799800 $Y=300460
X65 514 502 496 2 1 494 QDFFRBN $T=812820 315960 0 180 $X=801040 $Y=310540
X66 515 502 509 2 1 501 QDFFRBN $T=812820 326040 0 180 $X=801040 $Y=320620
X67 503 58 511 2 1 516 QDFFRBN $T=801040 346200 1 0 $X=801040 $Y=340780
X68 504 58 511 2 1 503 QDFFRBN $T=801040 346200 0 0 $X=801040 $Y=345820
X69 505 124 513 2 1 517 QDFFRBN $T=801040 356280 0 0 $X=801040 $Y=355900
X70 501 502 509 2 1 514 QDFFRBN $T=801660 315960 0 0 $X=801660 $Y=315580
X71 517 58 511 2 1 504 QDFFRBN $T=813440 356280 0 180 $X=801660 $Y=350860
X72 507 124 513 2 1 527 QDFFRBN $T=801660 366360 1 0 $X=801660 $Y=360940
X73 522 124 512 2 1 506 QDFFRBN $T=813440 386520 1 180 $X=801660 $Y=386140
X74 508 124 513 2 1 507 QDFFRBN $T=802280 366360 0 0 $X=802280 $Y=365980
X75 506 124 512 2 1 524 QDFFRBN $T=802280 386520 1 0 $X=802280 $Y=381100
X76 524 124 512 2 1 508 QDFFRBN $T=815300 376440 0 180 $X=803520 $Y=371020
X77 520 502 531 2 1 549 QDFFRBN $T=813440 305880 1 0 $X=813440 $Y=300460
X78 518 502 496 2 1 537 QDFFRBN $T=813440 305880 0 0 $X=813440 $Y=305500
X79 533 502 529 2 1 518 QDFFRBN $T=826460 315960 1 180 $X=814680 $Y=315580
X80 523 502 510 2 1 534 QDFFRBN $T=814680 336120 1 0 $X=814680 $Y=330700
X81 525 502 511 2 1 523 QDFFRBN $T=827080 346200 0 180 $X=815300 $Y=340780
X82 541 502 511 2 1 525 QDFFRBN $T=827080 346200 1 180 $X=815300 $Y=345820
X83 526 124 530 2 1 544 QDFFRBN $T=815300 366360 0 0 $X=815300 $Y=365980
X84 538 502 550 2 1 553 QDFFRBN $T=827080 315960 1 0 $X=827080 $Y=310540
X85 553 502 529 2 1 539 QDFFRBN $T=839480 326040 0 180 $X=827700 $Y=320620
X86 540 502 510 2 1 555 QDFFRBN $T=827700 336120 0 0 $X=827700 $Y=335740
X87 554 502 529 2 1 538 QDFFRBN $T=840100 305880 1 180 $X=828320 $Y=305500
X88 539 502 510 2 1 540 QDFFRBN $T=840100 336120 0 180 $X=828320 $Y=330700
X89 544 124 126 2 1 535 QDFFRBN $T=828320 366360 0 0 $X=828320 $Y=365980
X90 542 124 126 2 1 128 QDFFRBN $T=828320 386520 1 0 $X=828320 $Y=381100
X91 547 502 531 2 1 545 QDFFRBN $T=828940 295800 1 0 $X=828940 $Y=290380
X92 545 502 531 2 1 554 QDFFRBN $T=828940 295800 0 0 $X=828940 $Y=295420
X93 558 502 532 2 1 541 QDFFRBN $T=840720 346200 1 180 $X=828940 $Y=345820
X94 549 502 531 2 1 568 QDFFRBN $T=833900 305880 1 0 $X=833900 $Y=300460
X95 551 124 532 2 1 558 QDFFRBN $T=835760 366360 1 0 $X=835760 $Y=360940
X96 130 124 129 2 1 542 QDFFRBN $T=848160 386520 1 180 $X=836380 $Y=386140
X97 561 124 565 2 1 575 QDFFRBN $T=841960 356280 0 0 $X=841960 $Y=355900
X98 564 502 548 2 1 584 QDFFRBN $T=843820 275640 1 0 $X=843820 $Y=270220
X99 567 124 127 2 1 552 QDFFRBN $T=861180 376440 1 180 $X=849400 $Y=376060
X100 585 124 127 2 1 567 QDFFRBN $T=861180 386520 0 180 $X=849400 $Y=381100
X101 131 124 129 2 1 585 QDFFRBN $T=850020 386520 0 0 $X=850020 $Y=386140
X102 590 502 578 2 1 571 QDFFRBN $T=864280 305880 0 180 $X=852500 $Y=300460
X103 571 502 578 2 1 605 QDFFRBN $T=853740 295800 0 0 $X=853740 $Y=295420
X104 572 502 589 2 1 590 QDFFRBN $T=853740 315960 1 0 $X=853740 $Y=310540
X105 579 502 565 2 1 573 QDFFRBN $T=866760 336120 1 180 $X=854980 $Y=335740
X106 577 124 583 2 1 596 QDFFRBN $T=854980 366360 0 0 $X=854980 $Y=365980
X107 575 124 583 2 1 577 QDFFRBN $T=867380 356280 1 180 $X=855600 $Y=355900
X108 596 124 583 2 1 580 QDFFRBN $T=868000 376440 0 180 $X=856220 $Y=371020
X109 582 502 588 2 1 581 QDFFRBN $T=869240 285720 0 180 $X=857460 $Y=280300
X110 600 502 588 2 1 582 QDFFRBN $T=869860 275640 1 180 $X=858080 $Y=275260
X111 584 502 595 2 1 602 QDFFRBN $T=858700 275640 1 0 $X=858700 $Y=270220
X112 599 124 583 2 1 587 QDFFRBN $T=871720 356280 0 180 $X=859940 $Y=350860
X113 580 124 132 2 1 615 QDFFRBN $T=861800 386520 1 0 $X=861800 $Y=381100
X114 592 502 607 2 1 617 QDFFRBN $T=864280 305880 0 0 $X=864280 $Y=305500
X115 587 124 583 2 1 618 QDFFRBN $T=864280 366360 1 0 $X=864280 $Y=360940
X116 593 502 613 2 1 623 QDFFRBN $T=864900 336120 1 0 $X=864900 $Y=330700
X117 605 502 578 2 1 592 QDFFRBN $T=877300 305880 0 180 $X=865520 $Y=300460
X118 617 502 589 2 1 594 QDFFRBN $T=877300 326040 0 180 $X=865520 $Y=320620
X119 594 502 589 2 1 593 QDFFRBN $T=877300 326040 1 180 $X=865520 $Y=325660
X120 603 502 614 2 1 598 QDFFRBN $T=881640 336120 1 180 $X=869860 $Y=335740
X121 629 133 614 2 1 604 QDFFRBN $T=882260 356280 1 180 $X=870480 $Y=355900
X122 609 502 595 2 1 600 QDFFRBN $T=884120 275640 0 180 $X=872340 $Y=270220
X123 627 502 595 2 1 609 QDFFRBN $T=884120 275640 1 180 $X=872340 $Y=275260
X124 608 133 132 2 1 135 QDFFRBN $T=874820 386520 1 0 $X=874820 $Y=381100
X125 633 502 607 2 1 621 QDFFRBN $T=889080 315960 1 180 $X=877300 $Y=315580
X126 622 502 613 2 1 633 QDFFRBN $T=877920 326040 0 0 $X=877920 $Y=325660
X127 623 502 613 2 1 622 QDFFRBN $T=878540 336120 1 0 $X=878540 $Y=330700
X128 620 133 642 2 1 645 QDFFRBN $T=882880 366360 1 0 $X=882880 $Y=360940
X129 645 133 614 2 1 629 QDFFRBN $T=895280 356280 1 180 $X=883500 $Y=355900
X130 639 502 614 2 1 630 QDFFRBN $T=897760 336120 1 180 $X=885980 $Y=335740
X131 602 502 624 2 1 648 QDFFRBN $T=886600 275640 0 0 $X=886600 $Y=275260
X132 630 502 647 2 1 646 QDFFRBN $T=886600 346200 1 0 $X=886600 $Y=340780
X133 601 133 626 2 1 139 QDFFRBN $T=887220 386520 1 0 $X=887220 $Y=381100
X134 652 649 641 2 1 634 QDFFRBN $T=899620 295800 1 180 $X=887840 $Y=295420
X135 634 502 641 2 1 653 QDFFRBN $T=888460 305880 1 0 $X=888460 $Y=300460
X136 653 649 641 2 1 638 QDFFRBN $T=900860 305880 1 180 $X=889080 $Y=305500
X137 637 133 642 2 1 140 QDFFRBN $T=889080 366360 0 0 $X=889080 $Y=365980
X138 655 649 613 2 1 639 QDFFRBN $T=901480 326040 1 180 $X=889700 $Y=325660
X139 638 502 651 2 1 655 QDFFRBN $T=890320 315960 0 0 $X=890320 $Y=315580
X140 659 133 644 2 1 640 QDFFRBN $T=902100 376440 0 180 $X=890320 $Y=371020
X141 640 133 644 2 1 663 QDFFRBN $T=890940 376440 0 0 $X=890940 $Y=376060
X142 137 133 141 2 1 665 QDFFRBN $T=893420 386520 0 0 $X=893420 $Y=386140
X143 650 133 660 2 1 669 QDFFRBN $T=897760 356280 1 0 $X=897760 $Y=350860
X144 666 133 660 2 1 650 QDFFRBN $T=910160 356280 1 180 $X=898380 $Y=355900
X145 654 649 667 2 1 693 QDFFRBN $T=899620 265560 0 0 $X=899620 $Y=265180
X146 657 649 667 2 1 679 QDFFRBN $T=900240 275640 1 0 $X=900240 $Y=270220
X147 658 649 667 2 1 657 QDFFRBN $T=900240 275640 0 0 $X=900240 $Y=275260
X148 669 133 647 2 1 656 QDFFRBN $T=912020 346200 0 180 $X=900240 $Y=340780
X149 672 649 624 2 1 658 QDFFRBN $T=912640 285720 1 180 $X=900860 $Y=285340
X150 656 649 647 2 1 673 QDFFRBN $T=900860 336120 1 0 $X=900860 $Y=330700
X151 662 649 670 2 1 672 QDFFRBN $T=901480 295800 1 0 $X=901480 $Y=290380
X152 668 649 641 2 1 662 QDFFRBN $T=913880 305880 0 180 $X=902100 $Y=300460
X153 664 649 651 2 1 680 QDFFRBN $T=902100 315960 1 0 $X=902100 $Y=310540
X154 673 649 613 2 1 661 QDFFRBN $T=913880 326040 1 180 $X=902100 $Y=325660
X155 661 649 671 2 1 664 QDFFRBN $T=902720 326040 1 0 $X=902720 $Y=320620
X156 663 133 642 2 1 691 QDFFRBN $T=902720 366360 0 0 $X=902720 $Y=365980
X157 665 133 644 2 1 659 QDFFRBN $T=914500 376440 1 180 $X=902720 $Y=376060
X158 691 133 660 2 1 666 QDFFRBN $T=918220 366360 0 180 $X=906440 $Y=360940
X159 680 649 641 2 1 668 QDFFRBN $T=919460 305880 1 180 $X=907680 $Y=305500
X160 146 133 143 2 1 142 QDFFRBN $T=919460 386520 1 180 $X=907680 $Y=386140
X161 696 649 685 2 1 654 QDFFRBN $T=925040 265560 0 180 $X=913260 $Y=260140
X162 675 133 660 2 1 698 QDFFRBN $T=913260 346200 0 0 $X=913260 $Y=345820
X163 679 649 682 2 1 696 QDFFRBN $T=913880 275640 1 0 $X=913880 $Y=270220
X164 698 133 660 2 1 677 QDFFRBN $T=925660 356280 0 180 $X=913880 $Y=350860
X165 706 649 670 2 1 678 QDFFRBN $T=926280 285720 1 180 $X=914500 $Y=285340
X166 686 649 671 2 1 676 QDFFRBN $T=927520 326040 1 180 $X=915740 $Y=325660
X167 678 649 683 2 1 702 QDFFRBN $T=916360 295800 1 0 $X=916360 $Y=290380
X168 700 649 671 2 1 686 QDFFRBN $T=928140 326040 0 180 $X=916360 $Y=320620
X169 701 133 684 2 1 688 QDFFRBN $T=928140 376440 0 180 $X=916360 $Y=371020
X170 692 649 699 2 1 700 QDFFRBN $T=916980 315960 1 0 $X=916980 $Y=310540
X171 693 649 685 2 1 694 QDFFRBN $T=917600 265560 0 0 $X=917600 $Y=265180
X172 688 133 684 2 1 715 QDFFRBN $T=917600 366360 0 0 $X=917600 $Y=365980
X173 694 649 682 2 1 706 QDFFRBN $T=920080 275640 0 0 $X=920080 $Y=275260
X174 705 133 684 2 1 721 QDFFRBN $T=928140 376440 1 0 $X=928140 $Y=371020
X175 714 133 695 2 1 704 QDFFRBN $T=940540 336120 1 180 $X=928760 $Y=335740
X176 147 133 148 2 1 724 QDFFRBN $T=929380 386520 0 0 $X=929380 $Y=386140
X177 715 133 684 2 1 705 QDFFRBN $T=930000 366360 0 0 $X=930000 $Y=365980
X178 724 133 148 2 1 707 QDFFRBN $T=941780 386520 0 180 $X=930000 $Y=381100
X179 725 649 682 2 1 710 QDFFRBN $T=942400 275640 0 180 $X=930620 $Y=270220
X180 712 649 719 2 1 726 QDFFRBN $T=930620 295800 1 0 $X=930620 $Y=290380
X181 727 649 699 2 1 712 QDFFRBN $T=942400 305880 0 180 $X=930620 $Y=300460
X182 735 649 699 2 1 713 QDFFRBN $T=942400 305880 1 180 $X=930620 $Y=305500
X183 716 649 718 2 1 743 QDFFRBN $T=931240 245400 0 0 $X=931240 $Y=245020
X184 709 649 719 2 1 727 QDFFRBN $T=931240 315960 1 0 $X=931240 $Y=310540
X185 732 649 671 2 1 709 QDFFRBN $T=943020 336120 0 180 $X=931240 $Y=330700
X186 704 133 695 2 1 733 QDFFRBN $T=933100 346200 1 0 $X=933100 $Y=340780
X187 746 133 148 2 1 722 QDFFRBN $T=951700 376440 0 180 $X=939920 $Y=371020
X188 747 133 708 2 1 723 QDFFRBN $T=952320 356280 1 180 $X=940540 $Y=355900
X189 722 133 708 2 1 747 QDFFRBN $T=941160 366360 1 0 $X=941160 $Y=360940
X190 721 133 148 2 1 746 QDFFRBN $T=941160 376440 0 0 $X=941160 $Y=376060
X191 760 133 708 2 1 732 QDFFRBN $T=954180 336120 1 180 $X=942400 $Y=335740
X192 736 133 151 2 1 152 QDFFRBN $T=943640 386520 0 0 $X=943640 $Y=386140
X193 739 649 749 2 1 752 QDFFRBN $T=944260 285720 1 0 $X=944260 $Y=280300
X194 753 649 719 2 1 735 QDFFRBN $T=956040 305880 1 180 $X=944260 $Y=305500
X195 756 649 720 2 1 739 QDFFRBN $T=956660 275640 1 180 $X=944880 $Y=275260
X196 729 133 708 2 1 760 QDFFRBN $T=944880 346200 1 0 $X=944880 $Y=340780
X197 777 133 151 2 1 748 QDFFRBN $T=963480 376440 0 180 $X=951700 $Y=371020
X198 765 649 749 2 1 750 QDFFRBN $T=965340 285720 1 180 $X=953560 $Y=285340
X199 751 133 763 2 1 757 QDFFRBN $T=953560 346200 0 0 $X=953560 $Y=345820
X200 748 133 770 2 1 755 QDFFRBN $T=953560 366360 0 0 $X=953560 $Y=365980
X201 758 133 151 2 1 777 QDFFRBN $T=954800 376440 0 0 $X=954800 $Y=376060
X202 762 133 770 2 1 781 QDFFRBN $T=956660 346200 1 0 $X=956660 $Y=340780
X203 792 649 769 2 1 765 QDFFRBN $T=969680 295800 0 180 $X=957900 $Y=290380
X204 761 649 771 2 1 784 QDFFRBN $T=958520 315960 0 0 $X=958520 $Y=315580
X205 785 649 772 2 1 762 QDFFRBN $T=970300 336120 0 180 $X=958520 $Y=330700
X206 786 133 153 2 1 154 QDFFRBN $T=970300 386520 1 180 $X=958520 $Y=386140
X207 766 649 773 2 1 787 QDFFRBN $T=959140 275640 1 0 $X=959140 $Y=270220
X208 155 133 774 2 1 758 QDFFRBN $T=971540 386520 0 180 $X=959760 $Y=381100
X209 790 157 772 2 1 780 QDFFRBN $T=979600 336120 1 180 $X=967820 $Y=335740
X210 781 133 763 2 1 803 QDFFRBN $T=967820 346200 0 0 $X=967820 $Y=345820
X211 801 157 763 2 1 776 QDFFRBN $T=979600 356280 1 180 $X=967820 $Y=355900
X212 780 133 763 2 1 801 QDFFRBN $T=968440 346200 1 0 $X=968440 $Y=340780
X213 159 157 774 2 1 788 QDFFRBN $T=982080 386520 1 180 $X=970300 $Y=386140
X214 793 649 771 2 1 808 QDFFRBN $T=972160 326040 1 0 $X=972160 $Y=320620
X215 808 157 771 2 1 790 QDFFRBN $T=983940 336120 0 180 $X=972160 $Y=330700
X216 797 649 773 2 1 817 QDFFRBN $T=972780 265560 1 0 $X=972780 $Y=260140
X217 815 157 771 2 1 793 QDFFRBN $T=984560 315960 1 180 $X=972780 $Y=315580
X218 791 133 774 2 1 810 QDFFRBN $T=972780 366360 0 0 $X=972780 $Y=365980
X219 814 800 773 2 1 796 QDFFRBN $T=985180 265560 1 180 $X=973400 $Y=265180
X220 798 649 789 2 1 815 QDFFRBN $T=973400 305880 0 0 $X=973400 $Y=305500
X221 796 800 773 2 1 811 QDFFRBN $T=974020 275640 1 0 $X=974020 $Y=270220
X222 806 800 789 2 1 798 QDFFRBN $T=985800 295800 0 180 $X=974020 $Y=290380
X223 795 800 789 2 1 792 QDFFRBN $T=985800 295800 1 180 $X=974020 $Y=295420
X224 807 800 789 2 1 795 QDFFRBN $T=985800 305880 0 180 $X=974020 $Y=300460
X225 825 157 805 2 1 802 QDFFRBN $T=991380 336120 1 180 $X=979600 $Y=335740
X226 803 157 805 2 1 825 QDFFRBN $T=980220 346200 1 0 $X=980220 $Y=340780
X227 802 157 772 2 1 833 QDFFRBN $T=981460 326040 0 0 $X=981460 $Y=325660
X228 809 157 819 2 1 812 QDFFRBN $T=983940 356280 0 0 $X=983940 $Y=355900
X229 810 157 819 2 1 816 QDFFRBN $T=983940 376440 0 0 $X=983940 $Y=376060
X230 812 157 819 2 1 826 QDFFRBN $T=984560 356280 1 0 $X=984560 $Y=350860
X231 813 157 819 2 1 809 QDFFRBN $T=996340 366360 0 180 $X=984560 $Y=360940
X232 834 157 819 2 1 813 QDFFRBN $T=996960 366360 1 180 $X=985180 $Y=365980
X233 816 157 819 2 1 161 QDFFRBN $T=985800 386520 1 0 $X=985800 $Y=381100
X234 833 800 824 2 1 807 QDFFRBN $T=998200 326040 0 180 $X=986420 $Y=320620
X235 835 800 778 2 1 818 QDFFRBN $T=999440 285720 0 180 $X=987660 $Y=280300
X236 820 800 824 2 1 822 QDFFRBN $T=987660 315960 1 0 $X=987660 $Y=310540
X237 821 800 828 2 1 835 QDFFRBN $T=988280 295800 0 0 $X=988280 $Y=295420
X238 841 800 824 2 1 820 QDFFRBN $T=1000060 315960 1 180 $X=988280 $Y=315580
X239 826 157 805 2 1 842 QDFFRBN $T=989520 346200 0 0 $X=989520 $Y=345820
X240 827 157 830 2 1 841 QDFFRBN $T=990140 336120 1 0 $X=990140 $Y=330700
X241 842 157 830 2 1 827 QDFFRBN $T=1003160 336120 1 180 $X=991380 $Y=335740
X242 829 800 823 2 1 851 QDFFRBN $T=992000 275640 1 0 $X=992000 $Y=270220
X243 163 157 839 2 1 831 QDFFRBN $T=1007500 376440 1 180 $X=995720 $Y=376060
X244 831 157 839 2 1 854 QDFFRBN $T=996960 376440 1 0 $X=996960 $Y=371020
X245 854 157 839 2 1 834 QDFFRBN $T=1009980 366360 1 180 $X=998200 $Y=365980
X246 851 800 823 2 1 837 QDFFRBN $T=1010600 265560 1 180 $X=998820 $Y=265180
X247 869 157 805 2 1 838 QDFFRBN $T=1010600 356280 0 180 $X=998820 $Y=350860
X248 837 800 823 2 1 863 QDFFRBN $T=999440 265560 1 0 $X=999440 $Y=260140
X249 818 800 850 2 1 829 QDFFRBN $T=999440 285720 1 0 $X=999440 $Y=280300
X250 843 800 848 2 1 864 QDFFRBN $T=1001920 315960 0 0 $X=1001920 $Y=315580
X251 861 800 828 2 1 844 QDFFRBN $T=1014940 305880 0 180 $X=1003160 $Y=300460
X252 864 157 830 2 1 845 QDFFRBN $T=1014940 336120 0 180 $X=1003160 $Y=330700
X253 845 157 830 2 1 846 QDFFRBN $T=1014940 336120 1 180 $X=1003160 $Y=335740
X254 846 157 857 2 1 869 QDFFRBN $T=1003780 346200 0 0 $X=1003780 $Y=345820
X255 849 157 871 2 1 865 QDFFRBN $T=1007500 376440 0 0 $X=1007500 $Y=376060
X256 858 800 856 2 1 878 QDFFRBN $T=1012460 275640 1 0 $X=1012460 $Y=270220
X257 878 800 850 2 1 859 QDFFRBN $T=1024240 285720 0 180 $X=1012460 $Y=280300
X258 859 800 850 2 1 860 QDFFRBN $T=1024240 285720 1 180 $X=1012460 $Y=285340
X259 884 157 871 2 1 855 QDFFRBN $T=1024860 356280 1 180 $X=1013080 $Y=355900
X260 865 157 871 2 1 880 QDFFRBN $T=1013080 366360 0 0 $X=1013080 $Y=365980
X261 867 157 857 2 1 872 QDFFRBN $T=1013700 346200 1 0 $X=1013700 $Y=340780
X262 883 800 848 2 1 868 QDFFRBN $T=1026720 315960 1 180 $X=1014940 $Y=315580
X263 872 157 857 2 1 886 QDFFRBN $T=1014940 336120 0 0 $X=1014940 $Y=335740
X264 880 157 896 2 1 891 QDFFRBN $T=1023620 366360 1 0 $X=1023620 $Y=360940
X265 903 800 895 2 1 882 QDFFRBN $T=1037880 275640 1 180 $X=1026100 $Y=275260
X266 888 800 870 2 1 903 QDFFRBN $T=1026100 285720 0 0 $X=1026100 $Y=285340
X267 904 157 896 2 1 884 QDFFRBN $T=1037880 356280 1 180 $X=1026100 $Y=355900
X268 889 800 895 2 1 907 QDFFRBN $T=1026720 285720 1 0 $X=1026720 $Y=280300
X269 887 800 853 2 1 888 QDFFRBN $T=1038500 295800 1 180 $X=1026720 $Y=295420
X270 907 800 853 2 1 892 QDFFRBN $T=1039120 305880 0 180 $X=1027340 $Y=300460
X271 908 800 853 2 1 887 QDFFRBN $T=1039120 305880 1 180 $X=1027340 $Y=305500
X272 890 157 900 2 1 918 QDFFRBN $T=1027340 336120 1 0 $X=1027340 $Y=330700
X273 893 157 900 2 1 904 QDFFRBN $T=1027340 336120 0 0 $X=1027340 $Y=335740
X274 886 800 901 2 1 908 QDFFRBN $T=1027960 315960 0 0 $X=1027960 $Y=315580
X275 892 157 900 2 1 893 QDFFRBN $T=1027960 326040 0 0 $X=1027960 $Y=325660
X276 899 157 874 2 1 925 QDFFRBN $T=1036020 366360 0 0 $X=1036020 $Y=365980
X277 926 800 894 2 1 909 QDFFRBN $T=1050280 265560 0 180 $X=1038500 $Y=260140
X278 925 157 900 2 1 910 QDFFRBN $T=1050900 356280 1 180 $X=1039120 $Y=355900
X279 914 800 894 2 1 928 QDFFRBN $T=1039740 255480 0 0 $X=1039740 $Y=255100
X280 910 157 900 2 1 927 QDFFRBN $T=1039740 356280 1 0 $X=1039740 $Y=350860
X281 927 172 919 2 1 913 QDFFRBN $T=1052140 346200 0 180 $X=1040360 $Y=340780
X282 928 800 920 2 1 912 QDFFRBN $T=1052760 265560 1 180 $X=1040980 $Y=265180
X283 913 157 922 2 1 935 QDFFRBN $T=1040980 336120 0 0 $X=1040980 $Y=335740
X284 929 800 870 2 1 915 QDFFRBN $T=1053380 295800 1 180 $X=1041600 $Y=295420
X285 915 800 901 2 1 883 QDFFRBN $T=1053380 305880 1 180 $X=1041600 $Y=305500
X286 931 172 922 2 1 916 QDFFRBN $T=1053380 326040 0 180 $X=1041600 $Y=320620
X287 918 157 922 2 1 931 QDFFRBN $T=1041600 336120 1 0 $X=1041600 $Y=330700
X288 917 800 870 2 1 929 QDFFRBN $T=1042220 295800 1 0 $X=1042220 $Y=290380
X289 937 172 874 2 1 921 QDFFRBN $T=1057720 376440 0 180 $X=1045940 $Y=371020
X290 938 172 874 2 1 924 QDFFRBN $T=1058340 376440 1 180 $X=1046560 $Y=376060
X291 912 800 920 2 1 939 QDFFRBN $T=1047180 275640 1 0 $X=1047180 $Y=270220
X292 947 800 920 2 1 926 QDFFRBN $T=1062680 265560 0 180 $X=1050900 $Y=260140
X293 932 172 940 2 1 948 QDFFRBN $T=1051520 326040 0 0 $X=1051520 $Y=325660
X294 934 172 919 2 1 949 QDFFRBN $T=1052760 346200 0 0 $X=1052760 $Y=345820
X295 949 172 936 2 1 933 QDFFRBN $T=1064540 356280 1 180 $X=1052760 $Y=355900
X296 948 172 919 2 1 934 QDFFRBN $T=1065160 346200 0 180 $X=1053380 $Y=340780
X297 933 172 936 2 1 953 QDFFRBN $T=1053380 366360 1 0 $X=1053380 $Y=360940
X298 953 172 946 2 1 938 QDFFRBN $T=1069500 376440 0 180 $X=1057720 $Y=371020
X299 923 172 946 2 1 956 QDFFRBN $T=1059580 376440 0 0 $X=1059580 $Y=376060
X300 942 800 950 2 1 955 QDFFRBN $T=1060200 285720 0 0 $X=1060200 $Y=285340
X301 944 172 946 2 1 173 QDFFRBN $T=1060200 386520 0 0 $X=1060200 $Y=386140
X302 939 800 920 2 1 942 QDFFRBN $T=1072600 275640 0 180 $X=1060820 $Y=270220
X303 954 800 950 2 1 945 QDFFRBN $T=1072600 285720 0 180 $X=1060820 $Y=280300
X304 945 800 920 2 1 957 QDFFRBN $T=1061440 265560 0 0 $X=1061440 $Y=265180
X305 957 800 920 2 1 947 QDFFRBN $T=1074460 265560 0 180 $X=1062680 $Y=260140
X306 964 800 940 2 1 932 QDFFRBN $T=1075700 326040 1 180 $X=1063920 $Y=325660
X307 935 172 940 2 1 969 QDFFRBN $T=1065160 336120 0 0 $X=1065160 $Y=335740
X308 965 172 951 2 1 937 QDFFRBN $T=1077560 366360 1 180 $X=1065780 $Y=365980
X309 958 172 951 2 1 976 QDFFRBN $T=1073220 376440 1 0 $X=1073220 $Y=371020
X310 956 172 946 2 1 958 QDFFRBN $T=1085620 376440 1 180 $X=1073840 $Y=376060
X311 982 172 946 2 1 944 QDFFRBN $T=1085620 386520 1 180 $X=1073840 $Y=386140
X312 960 800 968 2 1 961 QDFFRBN $T=1075080 315960 1 0 $X=1075080 $Y=310540
X313 961 800 974 2 1 981 QDFFRBN $T=1075080 326040 1 0 $X=1075080 $Y=320620
X314 980 800 968 2 1 963 QDFFRBN $T=1087480 305880 1 180 $X=1075700 $Y=305500
X315 981 172 940 2 1 964 QDFFRBN $T=1088100 326040 1 180 $X=1076320 $Y=325660
X316 969 172 940 2 1 970 QDFFRBN $T=1078180 336120 0 0 $X=1078180 $Y=335740
X317 970 172 974 2 1 988 QDFFRBN $T=1079420 336120 1 0 $X=1079420 $Y=330700
X318 983 800 968 2 1 972 QDFFRBN $T=1092440 295800 0 180 $X=1080660 $Y=290380
X319 984 172 975 2 1 971 QDFFRBN $T=1093060 356280 0 180 $X=1081280 $Y=350860
X320 973 172 975 2 1 984 QDFFRBN $T=1081900 356280 0 0 $X=1081900 $Y=355900
X321 977 172 975 2 1 973 QDFFRBN $T=1094300 366360 0 180 $X=1082520 $Y=360940
X322 988 800 974 2 1 980 QDFFRBN $T=1099260 326040 0 180 $X=1087480 $Y=320620
X323 985 172 989 2 1 996 QDFFRBN $T=1092440 376440 0 0 $X=1092440 $Y=376060
X324 174 172 989 2 1 985 QDFFRBN $T=1104840 386520 0 180 $X=1093060 $Y=381100
X325 999 172 989 2 1 982 QDFFRBN $T=1105460 386520 1 180 $X=1093680 $Y=386140
X326 991 172 994 2 1 990 QDFFRBN $T=1096160 346200 1 0 $X=1096160 $Y=340780
X327 992 172 994 2 1 998 QDFFRBN $T=1096780 356280 0 0 $X=1096780 $Y=355900
X328 993 172 995 2 1 1002 QDFFRBN $T=1097400 366360 1 0 $X=1097400 $Y=360940
X329 996 172 995 2 1 992 QDFFRBN $T=1109180 376440 0 180 $X=1097400 $Y=371020
X330 1003 172 989 2 1 999 QDFFRBN $T=1120960 386520 1 180 $X=1109180 $Y=386140
X331 1000 172 989 2 1 1003 QDFFRBN $T=1109800 386520 1 0 $X=1109800 $Y=381100
X332 1002 172 995 2 1 1001 QDFFRBN $T=1110420 366360 1 0 $X=1110420 $Y=360940
X333 1001 172 995 2 1 1004 QDFFRBN $T=1110420 366360 0 0 $X=1110420 $Y=365980
X334 1004 172 989 2 1 1000 QDFFRBN $T=1122820 376440 1 180 $X=1111040 $Y=376060
X335 25 2 215 1 INV1S $T=553040 386520 0 180 $X=551800 $Y=381100
X336 26 2 217 1 INV1S $T=558000 376440 1 180 $X=556760 $Y=376060
X337 224 2 227 1 INV1S $T=561720 366360 0 0 $X=561720 $Y=365980
X338 232 2 239 1 INV1S $T=575360 366360 1 180 $X=574120 $Y=365980
X339 34 2 234 1 INV1S $T=577840 376440 1 0 $X=577840 $Y=371020
X340 211 2 249 1 INV1S $T=586520 376440 1 0 $X=586520 $Y=371020
X341 241 2 250 1 INV1S $T=587140 356280 1 0 $X=587140 $Y=350860
X342 257 2 273 1 INV1S $T=593340 376440 1 0 $X=593340 $Y=371020
X343 236 2 263 1 INV1S $T=596440 366360 0 0 $X=596440 $Y=365980
X344 253 2 265 1 INV1S $T=596440 376440 0 0 $X=596440 $Y=376060
X345 252 2 262 1 INV1S $T=597060 356280 0 0 $X=597060 $Y=355900
X346 40 2 269 1 INV1S $T=598920 386520 1 0 $X=598920 $Y=381100
X347 267 2 270 1 INV1S $T=600780 356280 1 0 $X=600780 $Y=350860
X348 272 2 264 1 INV1S $T=605740 366360 0 180 $X=604500 $Y=360940
X349 266 2 285 1 INV1S $T=613180 386520 1 180 $X=611940 $Y=386140
X350 258 2 288 1 INV1S $T=612560 356280 0 0 $X=612560 $Y=355900
X351 292 2 297 1 INV1S $T=620620 376440 0 0 $X=620620 $Y=376060
X352 311 2 318 1 INV1S $T=637980 376440 1 0 $X=637980 $Y=371020
X353 300 2 316 1 INV1S $T=639220 376440 0 0 $X=639220 $Y=376060
X354 62 2 322 1 INV1S $T=663400 376440 0 0 $X=663400 $Y=376060
X355 336 2 343 1 INV1S $T=680140 376440 1 0 $X=680140 $Y=371020
X356 338 2 347 1 INV1S $T=683240 376440 1 0 $X=683240 $Y=371020
X357 79 2 335 1 INV1S $T=684480 376440 0 0 $X=684480 $Y=376060
X358 84 2 357 1 INV1S $T=689440 386520 0 0 $X=689440 $Y=386140
X359 85 2 340 1 INV1S $T=690680 376440 0 0 $X=690680 $Y=376060
X360 83 2 361 1 INV1S $T=691300 366360 0 0 $X=691300 $Y=365980
X361 358 2 363 1 INV1S $T=692540 376440 0 0 $X=692540 $Y=376060
X362 372 2 364 1 INV1S $T=701840 376440 1 180 $X=700600 $Y=376060
X363 367 2 374 1 INV1S $T=701220 376440 1 0 $X=701220 $Y=371020
X364 375 2 380 1 INV1S $T=707420 386520 1 0 $X=707420 $Y=381100
X365 369 2 387 1 INV1S $T=712380 376440 0 0 $X=712380 $Y=376060
X366 366 2 396 1 INV1S $T=718580 356280 1 0 $X=718580 $Y=350860
X367 386 2 400 1 INV1S $T=720440 346200 1 0 $X=720440 $Y=340780
X368 98 2 401 1 INV1S $T=721060 386520 0 0 $X=721060 $Y=386140
X369 404 2 405 1 INV1S $T=724780 346200 1 0 $X=724780 $Y=340780
X370 101 2 412 1 INV1S $T=727260 386520 1 0 $X=727260 $Y=381100
X371 407 2 413 1 INV1S $T=729120 346200 0 0 $X=729120 $Y=345820
X372 408 2 420 1 INV1S $T=732220 376440 0 0 $X=732220 $Y=376060
X373 351 2 422 1 INV1S $T=732840 366360 1 0 $X=732840 $Y=360940
X374 419 2 421 1 INV1S $T=733460 346200 0 0 $X=733460 $Y=345820
X375 422 2 423 1 INV1S $T=734080 366360 1 0 $X=734080 $Y=360940
X376 433 2 430 1 INV1S $T=740280 376440 0 0 $X=740280 $Y=376060
X377 394 2 440 1 INV1S $T=743380 346200 1 0 $X=743380 $Y=340780
X378 435 2 458 1 INV1S $T=755780 356280 1 0 $X=755780 $Y=350860
X379 446 2 462 1 INV1S $T=757020 346200 1 0 $X=757020 $Y=340780
X380 425 2 468 1 INV1S $T=761360 356280 1 0 $X=761360 $Y=350860
X381 453 2 474 1 INV1S $T=764460 376440 1 0 $X=764460 $Y=371020
X382 467 2 475 1 INV1S $T=766320 386520 1 0 $X=766320 $Y=381100
X383 460 2 480 1 INV1S $T=767560 376440 0 0 $X=767560 $Y=376060
X384 535 2 576 1 INV1S $T=851260 376440 1 0 $X=851260 $Y=371020
X385 586 2 588 1 INV1S $T=859940 285720 0 0 $X=859940 $Y=285340
X386 567 2 597 1 INV1S $T=864280 376440 0 0 $X=864280 $Y=376060
X387 618 2 616 1 INV1S $T=876060 366360 1 180 $X=874820 $Y=365980
X388 615 2 611 1 INV1S $T=874820 376440 0 0 $X=874820 $Y=376060
X389 622 2 635 1 INV1S $T=889080 346200 0 0 $X=889080 $Y=345820
X390 646 2 643 1 INV1S $T=894040 346200 1 180 $X=892800 $Y=345820
X391 650 2 674 1 INV1S $T=909540 356280 1 0 $X=909540 $Y=350860
X392 677 2 687 1 INV1S $T=918840 356280 0 0 $X=918840 $Y=355900
X393 733 2 734 1 INV1S $T=943020 346200 0 0 $X=943020 $Y=345820
X394 729 2 744 1 INV1S $T=945500 346200 0 0 $X=945500 $Y=345820
X395 776 2 779 1 INV1S $T=965960 366360 1 0 $X=965960 $Y=360940
X396 803 2 794 1 INV1S $T=978980 356280 0 180 $X=977740 $Y=350860
X397 826 2 840 1 INV1S $T=998200 356280 0 0 $X=998200 $Y=355900
X398 838 2 847 1 INV1S $T=1003780 356280 0 0 $X=1003780 $Y=355900
X399 855 2 852 1 INV1S $T=1011220 356280 1 180 $X=1009980 $Y=355900
X400 872 2 866 1 INV1S $T=1018040 356280 0 180 $X=1016800 $Y=350860
X401 899 2 911 1 INV1S $T=1041600 386520 1 0 $X=1041600 $Y=381100
X402 924 2 902 1 INV1S $T=1047180 386520 0 180 $X=1045940 $Y=381100
X403 874 2 941 1 INV1S $T=1050900 366360 0 0 $X=1050900 $Y=365980
X404 941 2 951 1 INV1S $T=1062680 366360 0 0 $X=1062680 $Y=365980
X405 234 232 237 34 2 1 MXL2HS $T=569780 376440 0 0 $X=569780 $Y=376060
X406 404 450 455 405 2 1 MXL2HS $T=750200 346200 1 0 $X=750200 $Y=340780
X407 446 466 469 462 2 1 MXL2HS $T=760740 346200 1 0 $X=760740 $Y=340780
X408 419 476 483 421 2 1 MXL2HS $T=770040 346200 0 0 $X=770040 $Y=345820
X409 611 606 601 597 2 1 MXL2HS $T=873580 376440 1 180 $X=868000 $Y=376060
X410 616 606 608 576 2 1 MXL2HS $T=876060 376440 0 180 $X=870480 $Y=371020
X411 643 606 637 635 2 1 MXL2HS $T=892800 356280 0 180 $X=887220 $Y=350860
X412 687 606 144 674 2 1 MXL2HS $T=917600 356280 1 180 $X=912020 $Y=355900
X413 734 606 736 744 2 1 MXL2HS $T=942400 356280 1 0 $X=942400 $Y=350860
X414 779 606 786 794 2 1 MXL2HS $T=968440 366360 1 0 $X=968440 $Y=360940
X415 847 158 162 840 2 1 MXL2HS $T=1005640 366360 0 180 $X=1000060 $Y=360940
X416 852 158 165 866 2 1 MXL2HS $T=1009360 366360 1 0 $X=1009360 $Y=360940
X417 902 158 171 911 2 1 MXL2HS $T=1035400 386520 1 0 $X=1035400 $Y=381100
X418 138 502 1 2 INV12CK $T=895900 346200 0 0 $X=895900 $Y=345820
X419 138 649 1 2 INV12CK $T=932480 346200 0 0 $X=932480 $Y=345820
X420 156 133 1 2 INV12CK $T=975880 376440 0 180 $X=965960 $Y=371020
X421 156 800 1 2 INV12CK $T=982700 315960 0 180 $X=972780 $Y=310540
X422 156 157 1 2 INV12CK $T=996960 386520 1 180 $X=987040 $Y=386140
X423 250 242 1 2 267 AN2 $T=588380 356280 1 0 $X=588380 $Y=350860
X424 249 212 1 2 257 AN2 $T=589620 376440 1 0 $X=589620 $Y=371020
X425 400 392 1 2 404 AN2 $T=722300 346200 1 0 $X=722300 $Y=340780
X426 413 411 1 2 419 AN2 $T=730980 346200 0 0 $X=730980 $Y=345820
X427 478 480 1 2 485 AN2 $T=771900 376440 0 0 $X=771900 $Y=376060
X428 210 214 208 1 2 ND2 $T=549320 376440 0 180 $X=547460 $Y=371020
X429 210 222 221 1 2 ND2 $T=550560 376440 1 0 $X=550560 $Y=371020
X430 221 223 208 1 2 ND2 $T=554280 376440 1 0 $X=554280 $Y=371020
X431 218 236 229 1 2 ND2 $T=568540 376440 0 180 $X=566680 $Y=371020
X432 220 242 235 1 2 ND2 $T=579080 356280 1 180 $X=577220 $Y=355900
X433 38 246 37 1 2 ND2 $T=584040 386520 1 180 $X=582180 $Y=386140
X434 248 282 277 1 2 ND2 $T=608220 376440 1 180 $X=606360 $Y=376060
X435 281 286 287 1 2 ND2 $T=611320 366360 1 0 $X=611320 $Y=360940
X436 288 283 287 1 2 ND2 $T=614420 356280 0 0 $X=614420 $Y=355900
X437 287 298 262 1 2 ND2 $T=626200 356280 0 0 $X=626200 $Y=355900
X438 244 306 262 1 2 ND2 $T=631160 356280 1 180 $X=629300 $Y=355900
X439 316 315 294 1 2 ND2 $T=636740 376440 1 180 $X=634880 $Y=376060
X440 341 339 337 1 2 ND2 $T=679520 346200 1 180 $X=677660 $Y=345820
X441 342 337 345 1 2 ND2 $T=681380 346200 0 0 $X=681380 $Y=345820
X442 88 342 373 1 2 ND2 $T=705560 366360 1 180 $X=703700 $Y=365980
X443 89 373 91 1 2 ND2 $T=703700 376440 0 0 $X=703700 $Y=376060
X444 92 381 380 1 2 ND2 $T=709900 386520 1 0 $X=709900 $Y=381100
X445 348 392 321 1 2 ND2 $T=714860 346200 0 180 $X=713000 $Y=340780
X446 325 394 370 1 2 ND2 $T=717960 346200 0 180 $X=716100 $Y=340780
X447 388 411 393 1 2 ND2 $T=728500 346200 1 180 $X=726640 $Y=345820
X448 409 418 416 1 2 ND2 $T=734700 356280 0 180 $X=732840 $Y=350860
X449 447 457 445 1 2 ND2 $T=750200 376440 0 180 $X=748340 $Y=371020
X450 448 452 444 1 2 ND2 $T=753300 356280 0 180 $X=751440 $Y=350860
X451 442 465 443 1 2 ND2 $T=758880 376440 1 180 $X=757020 $Y=376060
X452 474 477 457 1 2 ND2 $T=768800 376440 0 180 $X=766940 $Y=371020
X453 468 479 418 1 2 ND2 $T=770040 356280 0 180 $X=768180 $Y=350860
X454 480 481 465 1 2 ND2 $T=771280 386520 0 180 $X=769420 $Y=381100
X455 19 16 1 17 2 209 OAI12HS $T=541260 386520 1 180 $X=537540 $Y=386140
X456 215 217 1 219 2 221 OAI12HS $T=548700 376440 0 0 $X=548700 $Y=376060
X457 25 26 1 27 2 219 OAI12HS $T=554900 386520 1 0 $X=554900 $Y=381100
X458 34 232 1 238 2 240 OAI12HS $T=576600 376440 0 180 $X=572880 $Y=371020
X459 234 239 1 240 2 243 OAI12HS $T=576600 366360 0 0 $X=576600 $Y=365980
X460 236 211 1 212 2 245 OAI12HS $T=585280 376440 0 180 $X=581560 $Y=371020
X461 40 253 1 247 2 274 OAI12HS $T=601400 386520 1 0 $X=601400 $Y=381100
X462 79 340 1 74 2 334 OAI12HS $T=683240 376440 1 180 $X=679520 $Y=376060
X463 345 342 1 350 2 341 OAI12HS $T=683240 356280 1 0 $X=683240 $Y=350860
X464 355 83 1 346 2 359 OAI12HS $T=688200 366360 1 0 $X=688200 $Y=360940
X465 361 71 1 359 2 350 OAI12HS $T=691920 366360 1 0 $X=691920 $Y=360940
X466 90 89 1 381 2 378 OAI12HS $T=706180 386520 0 0 $X=706180 $Y=386140
X467 394 386 1 392 2 410 OAI12HS $T=729740 346200 0 180 $X=726020 $Y=340780
X468 408 433 1 424 2 428 OAI12HS $T=738420 376440 1 180 $X=734700 $Y=376060
X469 420 430 1 428 2 445 OAI12HS $T=735940 376440 1 0 $X=735940 $Y=371020
X470 465 453 1 457 2 459 OAI12HS $T=761360 376440 0 180 $X=757640 $Y=371020
X471 460 467 1 465 2 471 OAI12HS $T=763840 376440 0 0 $X=763840 $Y=376060
X472 231 218 1 229 2 NR2T $T=569160 366360 1 180 $X=564200 $Y=365980
X473 291 307 1 309 2 NR2T $T=631160 366360 1 0 $X=631160 $Y=360940
X474 223 1 214 229 2 222 ND3 $T=556760 376440 1 0 $X=556760 $Y=371020
X475 291 1 281 284 2 290 ND3 $T=618140 366360 0 180 $X=615660 $Y=360940
X476 291 1 262 299 2 290 ND3 $T=621240 356280 0 0 $X=621240 $Y=355900
X477 291 1 255 293 2 48 ND3 $T=625580 366360 0 180 $X=623100 $Y=360940
X478 316 1 313 310 2 290 ND3 $T=640460 376440 1 0 $X=640460 $Y=371020
X479 454 1 452 450 2 449 ND3 $T=753300 346200 1 180 $X=750820 $Y=345820
X480 458 1 456 463 2 451 ND3 $T=756400 356280 0 0 $X=756400 $Y=355900
X481 418 1 470 476 2 472 ND3 $T=764460 346200 0 0 $X=764460 $Y=345820
X482 468 1 456 472 2 451 ND3 $T=766940 356280 1 180 $X=764460 $Y=355900
X483 206 14 208 2 1 XNR2HS $T=532580 376440 0 0 $X=532580 $Y=376060
X484 28 225 226 2 1 XNR2HS $T=559240 366360 1 0 $X=559240 $Y=360940
X485 27 228 225 2 1 XNR2HS $T=565440 376440 1 180 $X=559860 $Y=376060
X486 25 26 228 2 1 XNR2HS $T=559860 386520 1 0 $X=559860 $Y=381100
X487 224 226 230 2 1 XNR2HS $T=561720 356280 0 0 $X=561720 $Y=355900
X488 38 37 254 2 1 XNR2HS $T=586520 386520 0 0 $X=586520 $Y=386140
X489 40 253 261 2 1 XNR2HS $T=592100 386520 1 0 $X=592100 $Y=381100
X490 41 254 266 2 1 XNR2HS $T=595820 386520 0 0 $X=595820 $Y=386140
X491 43 266 42 2 1 XNR2HS $T=610700 386520 1 180 $X=605120 $Y=386140
X492 301 305 308 2 1 XNR2HS $T=628060 386520 1 0 $X=628060 $Y=381100
X493 63 64 324 2 1 XNR2HS $T=662780 386520 0 0 $X=662780 $Y=386140
X494 67 327 329 2 1 XNR2HS $T=667740 376440 1 0 $X=667740 $Y=371020
X495 63 61 330 2 1 XNR2HS $T=668360 386520 1 0 $X=668360 $Y=381100
X496 329 344 351 2 1 XNR2HS $T=682620 366360 1 0 $X=682620 $Y=360940
X497 346 356 360 2 1 XNR2HS $T=688200 356280 1 0 $X=688200 $Y=350860
X498 75 86 367 2 1 XNR2HS $T=693780 386520 1 0 $X=693780 $Y=381100
X499 80 86 369 2 1 XNR2HS $T=694400 376440 0 0 $X=694400 $Y=376060
X500 88 61 375 2 1 XNR2HS $T=699980 386520 1 0 $X=699980 $Y=381100
X501 88 64 90 2 1 XNR2HS $T=700600 386520 0 0 $X=700600 $Y=386140
X502 71 93 389 2 1 XNR2HS $T=710520 366360 1 0 $X=710520 $Y=360940
X503 94 64 372 2 1 XNR2HS $T=710520 386520 0 0 $X=710520 $Y=386140
X504 389 368 399 2 1 XNR2HS $T=717340 366360 1 0 $X=717340 $Y=360940
X505 371 398 408 2 1 XNR2HS $T=722300 376440 0 0 $X=722300 $Y=376060
X506 101 102 415 2 1 XNR2HS $T=727260 386520 0 0 $X=727260 $Y=386140
X507 378 403 429 2 1 XNR2HS $T=732840 386520 0 0 $X=732840 $Y=386140
X508 103 429 438 2 1 XNR2HS $T=738420 386520 0 0 $X=738420 $Y=386140
X509 408 433 439 2 1 XNR2HS $T=740280 386520 1 0 $X=740280 $Y=381100
X510 424 439 442 2 1 XNR2HS $T=748960 376440 1 180 $X=743380 $Y=376060
X511 306 314 54 1 2 XOR2H $T=637980 356280 0 0 $X=637980 $Y=355900
X512 315 319 57 1 2 XOR2H $T=643560 376440 0 0 $X=643560 $Y=376060
X513 28 2 233 225 1 NR2 $T=569160 366360 0 0 $X=569160 $Y=365980
X514 256 2 259 251 1 NR2 $T=594580 366360 1 0 $X=594580 $Y=360940
X515 357 2 365 77 1 NR2 $T=691920 386520 0 0 $X=691920 $Y=386140
X516 87 2 371 365 1 NR2 $T=696880 386520 1 180 $X=695020 $Y=386140
X517 355 2 377 368 1 NR2 $T=701840 366360 1 0 $X=701840 $Y=360940
X518 321 2 386 348 1 NR2 $T=711140 346200 0 180 $X=709280 $Y=340780
X519 96 2 390 97 1 NR2 $T=716720 386520 0 0 $X=716720 $Y=386140
X520 102 2 417 412 1 NR2 $T=730360 386520 1 0 $X=730360 $Y=381100
X521 427 2 436 434 1 NR2 $T=740280 346200 0 0 $X=740280 $Y=345820
X522 395 2 446 440 1 NR2 $T=745240 346200 1 0 $X=745240 $Y=340780
X523 20 2 207 1 211 NR2P $T=544980 376440 0 180 $X=541260 $Y=371020
X524 235 2 220 1 241 NR2P $T=578460 366360 0 180 $X=574740 $Y=360940
X525 243 2 230 1 252 NR2P $T=584660 366360 0 180 $X=580940 $Y=360940
X526 256 2 258 1 255 NR2P $T=593960 366360 0 180 $X=590240 $Y=360940
X527 245 2 259 1 260 NR2P $T=595820 366360 1 180 $X=592100 $Y=365980
X528 231 2 251 1 271 NR2P $T=603260 366360 1 180 $X=599540 $Y=365980
X529 263 2 231 1 272 NR2P $T=600780 366360 1 0 $X=600780 $Y=360940
X530 263 2 271 1 278 NR2P $T=607600 366360 1 180 $X=603880 $Y=365980
X531 231 2 258 1 281 NR2P $T=609460 366360 0 180 $X=605740 $Y=360940
X532 370 2 325 1 395 NR2P $T=718580 346200 1 180 $X=714860 $Y=345820
X533 393 2 388 1 407 NR2P $T=724780 346200 1 180 $X=721060 $Y=345820
X534 409 2 414 1 425 NR2P $T=732220 356280 0 0 $X=732220 $Y=355900
X535 410 2 436 1 426 NR2P $T=741520 346200 0 180 $X=737800 $Y=340780
X536 427 2 435 1 441 NR2P $T=744620 356280 0 180 $X=740900 $Y=350860
X537 395 2 435 1 448 NR2P $T=750200 356280 0 180 $X=746480 $Y=350860
X538 445 2 447 1 453 NR2P $T=748960 366360 0 0 $X=748960 $Y=365980
X539 443 2 442 1 460 NR2P $T=752680 376440 0 0 $X=752680 $Y=376060
X540 108 2 111 1 478 NR2P $T=773760 386520 1 180 $X=770040 $Y=386140
X541 225 28 1 233 235 227 2 MOAI1 $T=567920 366360 1 0 $X=567920 $Y=360940
X542 340 336 1 76 332 335 2 MOAI1 $T=679520 376440 0 180 $X=675180 $Y=371020
X543 364 340 1 363 368 82 2 MOAI1 $T=693160 376440 1 0 $X=693160 $Y=371020
X544 355 368 1 377 383 93 2 MOAI1 $T=704940 366360 1 0 $X=704940 $Y=360940
X545 92 367 1 89 385 387 2 MOAI1 $T=708660 376440 1 0 $X=708660 $Y=371020
X546 97 96 1 371 391 390 2 MOAI1 $T=718580 386520 0 180 $X=714240 $Y=381100
X547 99 98 1 82 402 372 2 MOAI1 $T=726020 386520 0 180 $X=721680 $Y=381100
X548 100 99 1 82 403 401 2 MOAI1 $T=726640 386520 1 180 $X=722300 $Y=386140
X549 230 1 243 244 2 ND2P $T=585280 356280 1 180 $X=581560 $Y=355900
X550 246 1 39 253 2 ND2P $T=586520 386520 1 0 $X=586520 $Y=381100
X551 295 1 289 294 2 ND2P $T=621240 386520 0 180 $X=617520 $Y=381100
X552 287 1 255 296 2 ND2P $T=618760 366360 1 0 $X=618760 $Y=360940
X553 441 1 444 437 2 ND2P $T=745240 356280 0 0 $X=745240 $Y=355900
X554 383 366 382 1 2 393 MAO222 $T=711760 356280 1 0 $X=711760 $Y=350860
X555 403 378 103 1 2 433 MAO222 $T=732840 386520 1 0 $X=732840 $Y=381100
X556 218 18 2 209 213 1 207 FA1 $T=549320 386520 0 180 $X=533820 $Y=381100
X557 210 24 2 22 21 1 213 FA1 $T=543120 386520 0 0 $X=543120 $Y=386140
X558 238 29 2 30 32 1 224 FA1 $T=575980 386520 1 180 $X=560480 $Y=386140
X559 247 35 2 33 36 1 232 FA1 $T=584660 386520 0 180 $X=569160 $Y=381100
X560 321 331 2 334 323 1 344 FA1 $T=663400 366360 1 0 $X=663400 $Y=360940
X561 325 339 2 326 320 1 348 FA1 $T=668360 346200 1 0 $X=668360 $Y=340780
X562 353 72 2 71 333 1 326 FA1 $T=684480 356280 1 180 $X=668980 $Y=355900
X563 366 376 2 352 360 1 384 FA1 $T=696260 356280 1 0 $X=696260 $Y=350860
X564 388 362 2 353 384 1 370 FA1 $T=714240 346200 1 180 $X=698740 $Y=345820
X565 406 95 2 385 391 1 382 FA1 $T=724160 366360 1 180 $X=708660 $Y=365980
X566 424 379 2 402 417 1 397 FA1 $T=734700 376440 0 180 $X=719200 $Y=371020
X567 447 397 2 399 406 1 409 FA1 $T=741520 366360 1 180 $X=726020 $Y=365980
X568 106 105 2 415 438 1 443 FA1 $T=761360 386520 1 180 $X=745860 $Y=386140
X569 291 290 2 287 1 314 AOI12HS $T=633020 356280 0 0 $X=633020 $Y=355900
X570 313 290 2 318 1 319 AOI12HS $T=642940 376440 1 0 $X=642940 $Y=371020
X571 456 451 2 444 1 484 AOI12HS $T=769420 356280 0 0 $X=769420 $Y=355900
X572 16 15 206 2 1 XOR2HS $T=536300 386520 1 180 $X=530720 $Y=386140
X573 210 216 220 2 1 XOR2HS $T=548700 366360 1 0 $X=548700 $Y=360940
X574 208 221 216 2 1 XOR2HS $T=554280 366360 1 180 $X=548700 $Y=365980
X575 74 75 336 2 1 XOR2HS $T=674560 386520 1 0 $X=674560 $Y=381100
X576 74 80 338 2 1 XOR2HS $T=686960 386520 0 180 $X=681380 $Y=381100
X577 74 61 358 2 1 XOR2HS $T=687580 386520 1 0 $X=687580 $Y=381100
X578 71 83 356 2 1 XOR2HS $T=688200 356280 0 0 $X=688200 $Y=355900
X579 350 354 362 2 1 XOR2HS $T=688820 346200 0 0 $X=688820 $Y=345820
X580 96 97 398 2 1 XOR2HS $T=716100 376440 0 0 $X=716100 $Y=376060
X581 479 484 486 2 1 XOR2HS $T=771900 356280 1 0 $X=771900 $Y=350860
X582 477 487 489 2 1 XOR2HS $T=775620 376440 1 0 $X=775620 $Y=371020
X583 481 488 490 2 1 XOR2HS $T=779340 386520 1 0 $X=779340 $Y=381100
X584 92 88 1 89 374 376 2 MOAI1S $T=707420 376440 0 180 $X=703700 $Y=371020
X585 369 92 1 89 375 379 2 MOAI1S $T=711140 376440 1 180 $X=707420 $Y=376060
X586 207 212 20 2 1 ND2S $T=544980 376440 1 180 $X=543120 $Y=376060
X587 297 301 282 2 1 ND2S $T=623100 376440 0 0 $X=623100 $Y=376060
X588 444 461 458 2 1 ND2S $T=758260 356280 1 0 $X=758260 $Y=350860
X589 444 470 468 2 1 ND2S $T=765700 356280 0 180 $X=763840 $Y=350860
X590 45 43 1 46 295 285 2 MOAI1H $T=614420 386520 0 0 $X=614420 $Y=386140
X591 338 340 1 343 345 82 2 MOAI1H $T=677040 366360 0 0 $X=677040 $Y=365980
X592 340 358 1 335 352 347 2 MOAI1H $T=692540 376440 0 180 $X=685100 $Y=371020
X593 273 276 1 2 INV2 $T=605120 376440 1 0 $X=605120 $Y=371020
X594 307 313 1 2 INV2 $T=634260 376440 1 0 $X=634260 $Y=371020
X595 51 317 1 2 INV2 $T=639840 386520 0 0 $X=639840 $Y=386140
X596 345 349 1 2 INV2 $T=684480 346200 0 0 $X=684480 $Y=345820
X597 71 355 1 2 INV2 $T=698740 366360 1 0 $X=698740 $Y=360940
X598 459 464 1 2 INV2 $T=758260 366360 0 0 $X=758260 $Y=365980
X599 478 482 1 2 INV2 $T=770040 376440 1 0 $X=770040 $Y=371020
X600 548 586 1 2 INV2 $T=849400 285720 0 0 $X=849400 $Y=285340
X601 586 595 1 2 INV2 $T=865520 285720 0 0 $X=865520 $Y=285340
X602 681 153 1 2 INV2 $T=957900 386520 0 180 $X=956040 $Y=381100
X603 681 769 1 2 INV2 $T=962240 295800 0 0 $X=962240 $Y=295420
X604 968 966 1 2 INV2 $T=1078800 295800 0 180 $X=1076940 $Y=290380
X605 966 967 1 2 INV2 $T=1080040 285720 0 0 $X=1080040 $Y=285340
X606 113 112 1 2 BUF2 $T=779340 386520 1 180 $X=776240 $Y=386140
X607 114 496 1 2 BUF2 $T=797320 315960 0 0 $X=797320 $Y=315580
X608 118 512 1 2 BUF2 $T=805380 376440 0 0 $X=805380 $Y=376060
X609 512 530 1 2 BUF2 $T=819640 376440 0 0 $X=819640 $Y=376060
X610 496 529 1 2 BUF2 $T=821500 315960 1 0 $X=821500 $Y=310540
X611 530 532 1 2 BUF2 $T=829560 366360 1 0 $X=829560 $Y=360940
X612 530 127 1 2 BUF2 $T=829560 376440 0 0 $X=829560 $Y=376060
X613 531 548 1 2 BUF2 $T=837000 285720 0 0 $X=837000 $Y=285340
X614 563 510 1 2 BUF2 $T=847540 336120 0 180 $X=844440 $Y=330700
X615 532 565 1 2 BUF2 $T=848780 356280 1 0 $X=848780 $Y=350860
X616 565 583 1 2 BUF2 $T=854360 356280 1 0 $X=854360 $Y=350860
X617 589 607 1 2 BUF2 $T=870480 315960 1 0 $X=870480 $Y=310540
X618 613 614 1 2 BUF2 $T=894660 336120 0 180 $X=891560 $Y=330700
X619 647 613 1 2 BUF2 $T=900240 336120 0 180 $X=897140 $Y=330700
X620 642 660 1 2 BUF2 $T=900240 366360 1 0 $X=900240 $Y=360940
X621 626 641 1 2 BUF2 $T=902100 305880 0 0 $X=902100 $Y=305500
X622 667 624 1 2 BUF2 $T=908300 285720 0 180 $X=905200 $Y=280300
X623 660 647 1 2 BUF2 $T=916360 346200 1 0 $X=916360 $Y=340780
X624 647 695 1 2 BUF2 $T=920080 346200 1 0 $X=920080 $Y=340780
X625 683 682 1 2 BUF2 $T=924420 285720 1 0 $X=924420 $Y=280300
X626 695 708 1 2 BUF2 $T=932480 346200 1 180 $X=929380 $Y=345820
X627 720 718 1 2 BUF2 $T=947980 255480 0 0 $X=947980 $Y=255100
X628 770 772 1 2 BUF2 $T=962240 336120 0 0 $X=962240 $Y=335740
X629 151 770 1 2 BUF2 $T=970920 366360 1 180 $X=967820 $Y=365980
X630 769 778 1 2 BUF2 $T=968440 285720 0 0 $X=968440 $Y=285340
X631 158 606 1 2 BUF2 $T=980220 366360 0 180 $X=977120 $Y=360940
X632 778 828 1 2 BUF2 $T=994480 285720 0 0 $X=994480 $Y=285340
X633 772 830 1 2 BUF2 $T=1001300 346200 1 0 $X=1001300 $Y=340780
X634 828 853 1 2 BUF2 $T=1005640 295800 0 0 $X=1005640 $Y=295420
X635 830 857 1 2 BUF2 $T=1007500 346200 1 0 $X=1007500 $Y=340780
X636 824 848 1 2 BUF2 $T=1008120 326040 0 0 $X=1008120 $Y=325660
X637 857 871 1 2 BUF2 $T=1023000 356280 0 180 $X=1019900 $Y=350860
X638 853 895 1 2 BUF2 $T=1039120 295800 1 0 $X=1039120 $Y=290380
X639 895 894 1 2 BUF2 $T=1040980 275640 0 0 $X=1040980 $Y=275260
X640 894 920 1 2 BUF2 $T=1046560 275640 0 0 $X=1046560 $Y=275260
X641 919 940 1 2 BUF2 $T=1060200 336120 0 0 $X=1060200 $Y=335740
X642 936 919 1 2 BUF2 $T=1069500 346200 1 180 $X=1066400 $Y=345820
X643 974 968 1 2 BUF2 $T=1090580 315960 1 180 $X=1087480 $Y=315580
X644 940 974 1 2 BUF2 $T=1091820 326040 0 0 $X=1091820 $Y=325660
X645 303 309 1 2 INV3 $T=629920 376440 1 0 $X=629920 $Y=371020
X646 681 626 1 2 INV3 $T=914500 386520 0 180 $X=912020 $Y=381100
X647 941 936 1 2 INV3 $T=1057100 366360 0 0 $X=1057100 $Y=365980
X648 966 950 1 2 INV3 $T=1078800 285720 1 180 $X=1076320 $Y=285340
X649 68 1 69 70 328 330 2 OAI22S $T=668980 386520 0 0 $X=668980 $Y=386140
X650 330 1 69 77 333 324 2 OAI22S $T=674560 386520 0 0 $X=674560 $Y=386140
X651 324 1 69 77 346 78 2 OAI22S $T=680140 386520 0 0 $X=680140 $Y=386140
X652 323 2 62 332 328 1 320 FA1S $T=672080 366360 1 180 $X=660300 $Y=365980
X653 327 2 322 65 73 1 331 FA1S $T=664640 376440 0 0 $X=664640 $Y=376060
X654 231 211 1 256 2 OR2T $T=584660 366360 0 0 $X=584660 $Y=365980
X655 50 49 1 307 2 OR2T $T=637980 386520 1 180 $X=631780 $Y=386140
X656 453 460 1 473 2 OR2T $T=761980 366360 0 0 $X=761980 $Y=365980
X657 490 58 118 123 1 2 QDFFRBP $T=786780 386520 1 0 $X=786780 $Y=381100
X658 113 1 451 2 BUF4CK $T=779960 366360 0 180 $X=775000 $Y=360940
X659 149 1 681 2 BUF4CK $T=943640 386520 1 0 $X=943640 $Y=381100
X660 280 275 283 251 1 2 ND3P $T=612560 356280 1 180 $X=607600 $Y=355900
X661 284 279 286 278 1 2 ND3P $T=614420 366360 1 180 $X=609460 $Y=365980
X662 290 280 288 291 1 2 ND3P $T=616280 356280 0 0 $X=616280 $Y=355900
X663 293 47 260 296 1 2 ND3P $T=616900 366360 0 0 $X=616900 $Y=365980
X664 299 302 298 244 1 2 ND3P $T=623100 356280 1 0 $X=623100 $Y=350860
X665 431 432 426 437 1 2 ND3P $T=737180 356280 0 0 $X=737180 $Y=355900
X666 451 449 448 456 1 2 ND3P $T=749580 356280 0 0 $X=749580 $Y=355900
X667 451 431 441 456 1 2 ND3P $T=749580 366360 1 0 $X=749580 $Y=360940
X668 463 466 461 434 1 2 ND3P $T=757640 346200 0 0 $X=757640 $Y=345820
X669 252 241 258 1 2 OR2P $T=590240 356280 0 0 $X=590240 $Y=355900
X670 395 386 427 1 2 OR2P $T=730980 346200 1 0 $X=730980 $Y=340780
X671 425 407 435 1 2 OR2P $T=736560 356280 1 0 $X=736560 $Y=350860
X672 277 2 1 248 292 NR2F $T=611940 376440 0 0 $X=611940 $Y=376060
X673 295 2 1 289 300 NR2F $T=621240 386520 1 0 $X=621240 $Y=381100
X674 292 2 1 300 303 NR2F $T=628680 376440 0 180 $X=621860 $Y=371020
X675 317 2 1 52 311 NR2F $T=639220 386520 1 0 $X=639220 $Y=381100
X676 482 2 1 473 456 NR2F $T=769420 366360 0 0 $X=769420 $Y=365980
X677 469 58 495 117 1005 1 2 DFFRBP $T=782440 346200 1 0 $X=782440 $Y=340780
X678 483 58 495 119 1006 1 2 DFFRBP $T=782440 346200 0 0 $X=782440 $Y=345820
X679 312 58 495 120 1007 1 2 DFFRBP $T=782440 356280 0 0 $X=782440 $Y=355900
X680 455 58 495 121 1008 1 2 DFFRBP $T=782440 366360 0 0 $X=782440 $Y=365980
X681 473 467 1 464 444 2 OAI12HP $T=768180 366360 0 180 $X=757640 $Y=360940
X682 311 300 1 294 305 310 2 OAI112HS $T=638600 386520 0 180 $X=634260 $Y=381100
X683 308 58 59 60 1 2 1009 DFFRBN $T=648520 386520 1 0 $X=648520 $Y=381100
X684 489 58 495 115 1 2 1010 DFFRBN $T=781820 376440 1 0 $X=781820 $Y=371020
X685 486 58 495 116 1 2 1011 DFFRBN $T=782440 356280 1 0 $X=782440 $Y=350860
X686 667 1 2 670 BUF1CK $T=912640 285720 1 0 $X=912640 $Y=280300
X687 695 1 2 671 BUF1CK $T=926900 336120 1 0 $X=926900 $Y=330700
X688 269 265 1 274 277 2 OAI12H $T=600160 376440 0 0 $X=600160 $Y=376060
X689 478 112 2 488 475 1 AOI12H $T=772520 386520 1 0 $X=772520 $Y=381100
X690 485 112 2 487 471 1 AOI12H $T=775620 376440 0 0 $X=775620 $Y=376060
X691 383 382 396 2 1 414 XNR3 $T=719820 356280 0 0 $X=719820 $Y=355900
X692 382 383 396 2 1 416 XNR3 $T=720440 356280 1 0 $X=720440 $Y=350860
X693 272 275 268 264 1 2 MXL2H $T=607600 356280 1 180 $X=598920 $Y=355900
X694 276 279 44 273 1 2 MXL2H $T=608840 376440 1 0 $X=608840 $Y=371020
X695 267 302 312 270 1 2 MXL2H $T=628680 356280 1 0 $X=628680 $Y=350860
X696 422 432 104 423 1 2 MXL2H $T=737180 366360 1 0 $X=737180 $Y=360940
X697 53 1 290 2 BUF6CK $T=641080 366360 1 0 $X=641080 $Y=360940
X698 237 248 238 1 2 XNR2H $T=580320 376440 0 0 $X=580320 $Y=376060
X699 261 289 247 1 2 XNR2H $T=608220 386520 1 0 $X=608220 $Y=381100
X700 342 354 349 1 2 XNR2H $T=694400 346200 0 180 $X=685720 $Y=340780
X701 241 244 242 251 1 2 OA12P $T=585900 356280 0 0 $X=585900 $Y=355900
X702 294 292 282 304 1 2 OA12P $T=626820 376440 0 0 $X=626820 $Y=376060
X703 407 418 411 434 1 2 OA12P $T=735320 346200 0 0 $X=735320 $Y=345820
X704 108 109 107 467 1 2 OA12P $T=766940 386520 1 180 $X=762600 $Y=386140
X705 309 311 1 304 287 2 OAI12HT $T=642320 366360 1 180 $X=627440 $Y=365980
X706 516 58 510 2 1 499 499 58 510 515 205 ICV_20 $T=801040 336120 1 0 $X=801040 $Y=330700
X707 537 502 528 2 1 519 519 502 528 547 205 ICV_20 $T=814060 295800 1 0 $X=814060 $Y=290380
X708 534 502 510 2 1 521 521 502 529 533 205 ICV_20 $T=814680 326040 1 0 $X=814680 $Y=320620
X709 536 124 512 2 1 522 125 124 126 536 205 ICV_20 $T=815300 386520 1 0 $X=815300 $Y=381100
X710 543 124 532 2 1 561 555 502 532 543 205 ICV_20 $T=840720 356280 0 180 $X=828940 $Y=350860
X711 552 124 127 2 1 566 566 124 127 551 205 ICV_20 $T=848160 376440 0 180 $X=836380 $Y=371020
X712 556 502 550 2 1 569 568 502 550 556 205 ICV_20 $T=851880 315960 0 180 $X=840100 $Y=310540
X713 557 502 563 2 1 570 569 502 563 557 205 ICV_20 $T=851880 326040 0 180 $X=840100 $Y=320620
X714 573 502 589 2 1 591 591 502 563 572 205 ICV_20 $T=864900 326040 0 180 $X=853120 $Y=320620
X715 574 502 583 2 1 599 598 502 565 579 205 ICV_20 $T=867380 346200 0 180 $X=855600 $Y=340780
X716 604 124 614 2 1 625 625 502 614 603 205 ICV_20 $T=882260 346200 0 180 $X=870480 $Y=340780
X717 628 502 595 2 1 610 610 502 624 627 205 ICV_20 $T=872340 285720 1 0 $X=872340 $Y=280300
X718 619 502 595 2 1 612 612 502 595 628 205 ICV_20 $T=872960 295800 1 0 $X=872960 $Y=290380
X719 134 133 626 2 1 636 636 133 626 620 205 ICV_20 $T=889700 376440 0 180 $X=877920 $Y=371020
X720 632 502 624 2 1 652 648 502 624 632 205 ICV_20 $T=899000 285720 0 180 $X=887220 $Y=280300
X721 697 649 647 2 1 675 676 649 695 697 205 ICV_20 $T=913260 336120 1 0 $X=913260 $Y=330700
X722 723 133 708 2 1 703 703 133 695 729 205 ICV_20 $T=927520 356280 1 0 $X=927520 $Y=350860
X723 726 649 683 2 1 711 711 649 682 725 205 ICV_20 $T=930620 285720 1 0 $X=930620 $Y=280300
X724 728 649 671 2 1 714 713 649 671 728 205 ICV_20 $T=930620 326040 1 0 $X=930620 $Y=320620
X725 717 649 718 2 1 730 730 649 718 716 205 ICV_20 $T=943020 255480 0 180 $X=931240 $Y=250060
X726 710 649 720 2 1 731 731 649 718 717 205 ICV_20 $T=943020 265560 0 180 $X=931240 $Y=260140
X727 737 649 745 2 1 753 752 649 745 737 205 ICV_20 $T=956040 295800 0 180 $X=944260 $Y=290380
X728 742 649 749 2 1 756 741 649 720 742 205 ICV_20 $T=957280 265560 0 180 $X=945500 $Y=260140
X729 755 133 770 2 1 775 775 133 763 751 205 ICV_20 $T=965960 356280 0 180 $X=954180 $Y=350860
X730 767 649 771 2 1 785 784 649 771 767 205 ICV_20 $T=970300 326040 0 180 $X=958520 $Y=320620
X731 787 649 773 2 1 768 768 649 773 797 205 ICV_20 $T=959140 265560 1 0 $X=959140 $Y=260140
X732 799 649 778 2 1 806 811 800 778 799 205 ICV_20 $T=986420 285720 0 180 $X=974640 $Y=280300
X733 832 800 823 2 1 814 817 800 823 832 205 ICV_20 $T=985800 265560 1 0 $X=985800 $Y=260140
X734 822 800 828 2 1 836 836 800 828 821 205 ICV_20 $T=1000060 305880 0 180 $X=988280 $Y=300460
X735 164 157 166 2 1 873 873 157 839 849 205 ICV_20 $T=1018660 386520 0 180 $X=1006880 $Y=381100
X736 877 800 856 2 1 858 863 800 856 877 205 ICV_20 $T=1012460 265560 1 0 $X=1012460 $Y=260140
X737 879 800 870 2 1 861 860 800 870 879 205 ICV_20 $T=1012460 295800 1 0 $X=1012460 $Y=290380
X738 881 157 848 2 1 867 868 800 848 881 205 ICV_20 $T=1014320 326040 1 0 $X=1014320 $Y=320620
X739 170 157 169 2 1 875 875 157 169 897 205 ICV_20 $T=1021140 386520 1 0 $X=1021140 $Y=381100
X740 897 157 871 2 1 876 876 157 871 898 205 ICV_20 $T=1021760 376440 1 0 $X=1021760 $Y=371020
X741 891 157 900 2 1 906 906 157 857 890 205 ICV_20 $T=1038500 346200 0 180 $X=1026720 $Y=340780
X742 898 157 874 2 1 923 921 157 874 899 205 ICV_20 $T=1045940 376440 0 180 $X=1034160 $Y=371020
X743 916 800 922 2 1 930 930 800 901 917 205 ICV_20 $T=1053380 315960 0 180 $X=1041600 $Y=310540
X744 943 800 950 2 1 954 955 800 950 943 205 ICV_20 $T=1071980 295800 0 180 $X=1060200 $Y=290380
X745 952 172 936 2 1 965 971 172 936 952 205 ICV_20 $T=1078180 356280 0 180 $X=1066400 $Y=350860
X746 990 172 994 2 1 997 997 172 974 986 205 ICV_20 $T=1107940 336120 0 180 $X=1096160 $Y=330700
X747 149 874 1 2 INV2CK $T=1019280 376440 0 0 $X=1019280 $Y=376060
X748 497 58 114 2 1 492 491 58 114 497 205 ICV_22 $T=795460 326040 1 180 $X=783680 $Y=325660
X749 535 124 530 2 1 505 527 124 530 526 205 ICV_22 $T=827080 356280 1 180 $X=815300 $Y=355900
X750 560 502 548 2 1 546 546 502 548 562 205 ICV_22 $T=841340 275640 1 180 $X=829560 $Y=275260
X751 570 502 565 2 1 559 559 502 565 574 205 ICV_22 $T=853120 336120 1 180 $X=841340 $Y=335740
X752 562 502 548 2 1 564 581 502 548 560 205 ICV_22 $T=843200 275640 0 0 $X=843200 $Y=275260
X753 631 502 607 2 1 619 621 502 607 631 205 ICV_22 $T=888460 305880 1 180 $X=876680 $Y=305500
X754 702 649 683 2 1 689 689 649 699 692 205 ICV_22 $T=928760 295800 1 180 $X=916980 $Y=295420
X755 690 133 684 2 1 701 707 133 143 690 205 ICV_22 $T=917600 376440 0 0 $X=917600 $Y=376060
X756 738 649 745 2 1 764 754 649 719 738 205 ICV_22 $T=944260 315960 0 0 $X=944260 $Y=315580
X757 740 649 719 2 1 754 757 133 708 740 205 ICV_22 $T=944880 326040 0 0 $X=944880 $Y=325660
X758 743 649 718 2 1 759 759 649 718 741 205 ICV_22 $T=945500 245400 0 0 $X=945500 $Y=245020
X759 782 649 745 2 1 761 764 649 745 782 205 ICV_22 $T=969680 305880 1 180 $X=957900 $Y=305500
X760 783 649 769 2 1 766 750 649 778 783 205 ICV_22 $T=970300 275640 1 180 $X=958520 $Y=275260
X761 804 157 774 2 1 791 788 133 774 804 205 ICV_22 $T=983940 376440 1 180 $X=972160 $Y=376060
X762 844 800 853 2 1 862 862 800 848 843 205 ICV_22 $T=1002540 305880 0 0 $X=1002540 $Y=305500
X763 882 800 894 2 1 914 909 800 894 885 205 ICV_22 $T=1026100 255480 0 0 $X=1026100 $Y=255100
X764 885 800 894 2 1 905 905 800 895 889 205 ICV_22 $T=1026720 265560 0 0 $X=1026720 $Y=265180
X765 978 800 950 2 1 962 959 800 967 978 205 ICV_22 $T=1087480 265560 1 180 $X=1075700 $Y=265180
X766 962 800 967 2 1 983 979 800 967 959 205 ICV_22 $T=1075700 275640 0 0 $X=1075700 $Y=275260
X767 963 800 968 2 1 979 972 800 968 960 205 ICV_22 $T=1075700 295800 0 0 $X=1075700 $Y=295420
X768 987 172 975 2 1 977 976 172 975 987 205 ICV_22 $T=1096780 366360 1 180 $X=1085000 $Y=365980
X769 998 172 994 2 1 991 986 172 994 993 205 ICV_22 $T=1108560 346200 1 180 $X=1096780 $Y=345820
X770 268 58 118 122 1 2 1012 DFFRBT $T=786160 376440 0 0 $X=786160 $Y=376060
X771 167 2 1 TIE1 $T=1009980 225240 1 0 $X=1009980 $Y=219820
X772 395 434 394 2 1 454 OA12S $T=745240 346200 0 0 $X=745240 $Y=345820
.ENDS
***************************************
.SUBCKT ICV_26 1 2 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26
+ 27 28 49
** N=68 EP=23 IP=52 FDC=0
X0 11 2 2 2 12 2 13 YA2GSD $T=417140 0 0 0 $X=419990 $Y=0
X1 14 9 9 9 15 9 13 YA2GSD $T=756770 0 0 0 $X=759620 $Y=0
X2 16 9 10 10 17 10 13 YA2GSD $T=869980 0 0 0 $X=872830 $Y=0
X3 18 10 10 19 20 19 21 YA2GSD $T=983190 0 0 0 $X=986040 $Y=0
X4 22 19 19 19 23 24 21 YA2GSD $T=1096400 0 0 0 $X=1099250 $Y=0
X5 25 1 1 1 26 XMD $T=190720 0 0 0 $X=193570 $Y=0
X6 27 1 1 2 28 XMD $T=303930 0 0 0 $X=306780 $Y=0
.ENDS
***************************************
.SUBCKT ICV_27
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_28 1 2 3 4 5 6
** N=7 EP=6 IP=8 FDC=0
X0 3 2 2 4 5 4 1 YA2GSD $T=0 1146820 0 270 $X=0 $Y=1087050
.ENDS
***************************************
.SUBCKT ICV_29 1 2 3 4
** N=5 EP=4 IP=6 FDC=0
X0 1 2 2 2 3 XMD $T=0 1020980 0 270 $X=0 $Y=961210
.ENDS
***************************************
.SUBCKT ICV_30 2 3 4 10
** N=11 EP=4 IP=6 FDC=0
X0 3 2 2 2 4 XMD $T=0 895140 0 270 $X=0 $Y=835370
.ENDS
***************************************
.SUBCKT ICV_31
** N=13 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_32 1 2 3 4
** N=5 EP=4 IP=6 FDC=0
X0 3 2 2 2 1 XMD $T=0 517640 0 270 $X=0 $Y=457870
.ENDS
***************************************
.SUBCKT ICV_33 1 2 3 4 5 6
** N=8 EP=6 IP=12 FDC=0
X0 3 1 1 1 4 XMD $T=0 265960 0 270 $X=0 $Y=206190
X1 5 1 1 1 2 XMD $T=0 391800 0 270 $X=0 $Y=332030
.ENDS
***************************************
.SUBCKT ICV_34
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT CHIP o_data[7] o_data[11] o_data[10] o_data[6] o_data[5] o_data[3] o_data[4] clk rst_n layer_num[0] layer_num[1] i_data[0] o_data[12] o_data[13] VCC GND i_data[6] i_data[7] o_data[0] o_data[1]
+ o_data[2] o_data[8] o_data[9] o_data[14] i_data[5] i_data[4] i_data[3] i_data[1] i_data[2]
** N=1222 EP=29 IP=2540 FDC=0
X0 o_data[7] 64 1 8 1222 ICV_1 $T=1349740 870270 0 90 $X=1210240 $Y=873120
X2 o_data[11] 65 116 8 1222 ICV_3 $T=0 0 0 0 $X=1210200 $Y=1077400
X3 4 5 o_data[10] 8 1222 ICV_4 $T=0 0 0 0 $X=1210200 $Y=900200
X4 7 8 o_data[6] 511 1222 ICV_5 $T=0 0 0 0 $X=1210200 $Y=719600
X6 o_data[5] 67 871 857 1222 ICV_7 $T=0 0 0 0 $X=1210200 $Y=391200
X7 12 o_data[3] 68 857 o_data[4] 69 844 1222 ICV_8 $T=0 0 0 0 $X=1210200 $Y=139500
X9 16 25 28 30 o_data[12] 80 8 o_data[13] 81 clk 33 872 rst_n 70 layer_num[0] 77 layer_num[1] 78 i_data[0] 79
+ 1222
+ ICV_10 $T=0 0 0 0 $X=139500 $Y=1210660
X10 33 GND VCC 872 896 82 16 70 83 85 84 897 86 87 88 89 90 91 92 95
+ 93 97 94 96 98 898 99 899 100 101 25 102 103 104 105 106 107 112 108 109
+ 111 110 900 113 114 115 28 30 65 1222
+ ICV_11 $T=0 0 0 0 $X=139500 $Y=1076620
X11 GND VCC 36 82 121 127 118 117 119 120 125 83 122 902 123 942 124 901 224 903
+ 126 905 128 129 132 130 131 137 133 134 135 136 138 140 141 142 139 143 145 146
+ 144 84 912 154 904 897 147 149 162 148 85 86 152 906 150 907 151 153 155 156
+ 157 158 97 159 160 161 163 164 167 169 165 166 87 193 908 88 168 89 90 91
+ 170 179 909 172 92 171 93 174 175 173 95 94 176 177 911 178 96 913 180 181
+ 182 898 183 184 185 915 914 186 98 187 188 99 189 100 190 101 917 191 192 102
+ 899 195 194 196 916 103 198 197 104 106 105 918 199 204 200 919 201 202 203 206
+ 205 924 921 219 207 107 900 208 78 209 77 210 910 108 920 212 211 922 109 213
+ 110 214 215 111 112 216 113 218 114 217 220 221 881 115 222 225 925 223 926 927
+ 923 226 228 227 229 930 230 928 232 929 231 931 238 233 236 234 235 237 940 239
+ 240 952 241 243 242 256 244 245 248 936 246 937 947 948 262 247 932 249 250 252
+ 934 933 935 251 253 255 254 938 939 941 257 945 943 258 946 259 944 260 882 949
+ 883 950 275 951 263 261 264 265 954 953 266 267 956 884 268 269 957 960 955 270
+ 958 272 959 271 274 273 276 277 278 279 281 282 284 280 283 287 285 286 288 4
+ 64 65 1222
+ ICV_16 $T=0 0 0 0 $X=139500 $Y=900200
X12 GND VCC 289 290 291 293 962 292 961 295 294 298 296 297 299 963 300 301 302 303
+ 305 304 306 117 307 127 118 119 313 311 121 120 308 122 964 318 977 123 309 310
+ 125 124 312 901 323 903 314 315 965 967 316 317 126 968 969 319 320 970 972 321
+ 973 326 128 129 974 322 971 966 975 131 325 324 130 327 132 133 137 328 976 329
+ 134 330 336 331 332 140 333 334 979 978 335 135 136 980 138 142 337 981 139 338
+ 141 146 904 144 339 143 999 340 145 341 1002 902 342 985 983 982 984 367 993 343
+ 344 345 986 987 348 346 347 988 162 989 154 366 990 1003 349 350 351 147 352 991
+ 353 148 992 149 354 994 995 358 355 357 150 356 151 906 152 359 996 998 997 360
+ 153 1001 361 363 362 364 155 156 157 365 160 368 158 159 369 1007 370 371 372 1004
+ 373 374 161 165 375 1005 163 377 376 380 404 1000 164 166 379 167 193 908 378 1006
+ 381 169 399 170 383 384 382 1008 219 909 385 1009 386 910 168 171 172 173 920 174
+ 387 1010 1011 176 388 175 389 911 1012 177 178 390 912 391 1013 392 913 179 180 393
+ 181 182 394 183 184 395 396 1015 397 401 185 914 398 187 188 400 190 186 189 403
+ 402 192 916 1016 191 917 194 915 198 405 195 1014 196 406 197 921 407 408 413 409
+ 203 411 199 200 918 412 1021 416 1020 410 919 201 202 414 428 415 1018 1022 208 204
+ 1023 1024 417 423 205 206 212 418 1026 1032 1028 1027 419 420 207 1029 1030 210 1033 1031
+ 421 422 437 922 1037 424 209 1034 1035 211 1039 425 1036 426 427 436 213 881 214 429
+ 1038 1040 433 216 430 215 431 217 221 227 432 240 218 434 222 220 923 435 1049 438
+ 925 223 224 924 225 926 443 226 927 229 228 499 230 439 1043 930 440 929 233 1042
+ 928 231 232 441 237 235 238 234 931 442 239 236 455 1044 444 448 249 445 244 1041
+ 446 447 1045 1019 1046 242 449 1047 248 243 450 934 245 1017 241 247 246 1048 451 932
+ 454 452 933 453 268 250 251 936 253 456 935 255 252 254 457 937 948 938 1050 939
+ 884 941 256 458 460 940 261 459 258 259 1025 943 262 1051 945 1052 260 944 946 953
+ 462 882 947 461 1054 463 952 1055 265 464 1053 956 465 883 263 466 955 1056 954 1058
+ 950 264 467 468 266 470 267 469 269 471 1060 951 957 1059 958 472 271 959 474 272
+ 475 1061 949 473 276 273 1065 476 1057 1063 478 477 1064 960 275 274 479 1066 277 1068
+ 1062 480 481 270 485 482 279 278 483 1070 1069 484 282 280 1067 281 1071 283 486 942
+ 487 1072 286 284 285 489 490 501 287 491 288 488 492 493 495 506 494 496 497 498
+ 500 502 503 504 505 509 507 508 510 7 64 1222
+ ICV_19 $T=0 0 0 0 $X=139500 $Y=718780
X13 GND VCC 1078 512 513 514 290 517 1073 516 291 961 518 515 292 519 1074 520 962 293
+ 521 522 296 294 523 295 524 1075 1077 299 527 533 297 525 526 1076 298 528 963 530
+ 529 300 531 301 532 302 1079 303 534 978 304 305 536 306 537 535 539 540 538 309
+ 543 541 308 542 964 311 966 544 310 313 314 545 316 965 315 885 307 319 546 972
+ 318 547 971 880 317 321 548 968 969 1080 970 320 1082 550 549 553 1081 323 551 974
+ 973 322 552 975 976 324 312 979 554 325 967 326 328 977 327 557 329 330 555 1083
+ 332 336 331 556 333 980 1085 335 1084 337 338 334 1088 558 560 340 1086 559 1089 339
+ 341 1087 561 1090 981 1091 342 562 343 563 344 366 983 984 345 985 986 987 347 346
+ 903 989 988 348 574 835 565 990 349 567 350 566 351 1096 352 991 1095 992 1097 569
+ 994 1094 571 907 353 575 570 1092 905 354 572 355 564 356 357 576 358 579 1098 998
+ 982 996 573 1100 1093 1101 580 359 1099 360 578 1000 1102 362 1103 583 361 1105 363 365
+ 1106 1108 993 997 1104 1001 364 1002 581 1111 577 1113 1110 582 999 1114 584 79 1003 367
+ 585 1109 369 587 1107 1116 586 1115 1112 589 995 1117 1118 368 371 372 588 370 1119 591
+ 379 568 373 592 374 1005 593 375 1006 1121 404 376 594 377 1122 378 384 380 595 598
+ 767 1126 896 381 599 596 1123 590 382 1124 1008 1007 383 386 219 1010 1127 1125 385 602
+ 600 1128 1012 1130 601 1129 387 1011 605 388 389 392 390 391 1133 603 597 393 394 1134
+ 604 1013 1136 1132 1131 395 606 607 398 396 1015 1135 397 608 609 610 399 400 401 611
+ 1138 402 612 1120 1137 613 409 1139 1141 1041 405 1017 615 1025 1019 614 406 1009 616 407
+ 618 617 619 620 1018 408 417 1140 410 1021 1020 411 1033 1022 621 1032 413 622 414 624
+ 412 428 623 1024 415 625 421 1023 1027 416 1040 1031 627 418 626 1026 419 420 1028 1029
+ 424 1036 628 1030 422 423 1034 425 426 427 630 1037 631 636 1035 632 429 431 1038 633
+ 634 430 635 1039 432 637 433 434 641 638 642 435 437 436 640 438 643 1142 651 644
+ 439 645 646 639 1144 647 1145 648 441 1143 440 629 442 1148 443 1042 649 444 447 650
+ 445 1045 446 1147 1049 1146 652 448 654 1149 450 655 451 1150 1044 449 656 1046 1047 659
+ 657 1048 653 452 660 661 454 658 1151 455 456 1153 453 1152 1154 1155 1050 662 1156 663
+ 675 457 1157 664 666 665 1159 1158 673 458 667 668 670 459 460 669 1160 1161 1051 671
+ 672 461 1171 1052 1054 1053 1164 1162 462 463 1055 1163 674 466 1058 676 464 465 677 1059
+ 1056 1173 678 1166 1167 679 680 1057 467 1165 682 697 681 468 683 471 684 1061 469 1169
+ 1168 1170 470 685 1062 1060 472 473 686 474 475 1065 687 1063 476 478 477 1064 879 688
+ 689 1066 690 1070 708 479 1043 1067 691 480 481 482 1069 485 1068 693 692 483 1071 501
+ 694 484 1072 487 1172 695 486 696 488 698 489 490 699 491 700 493 492 496 701 81
+ 494 702 495 506 1174 497 80 703 498 116 713 704 499 500 1175 5 706 709 705 707
+ 504 502 503 710 505 711 507 712 508 725 714 715 509 510 716 718 717 722 719 721
+ 720 723 724 1222
+ ICV_21 $T=0 0 0 0 $X=139500 $Y=542380
X14 GND VCC 37 512 513 289 1078 515 514 1073 516 517 518 1074 519 520 525 521 522 523
+ 524 1147 1077 1075 526 527 1076 528 529 530 531 532 534 533 535 536 537 538 539 540
+ 541 542 543 547 544 545 546 548 549 550 1081 551 1082 552 1080 726 553 554 727 734
+ 555 1083 556 559 557 1084 728 562 732 729 1085 558 39 1087 1088 1086 560 730 731 965
+ 561 1090 1089 733 563 1091 564 1092 1093 1094 565 1105 566 1098 1004 1107 567 1095 1096 568
+ 1097 1099 569 578 570 1100 571 1101 575 585 574 572 573 735 576 1000 1102 1108 1112 1103
+ 1104 577 1106 1121 1110 579 738 580 736 739 1113 581 1119 737 1114 582 1109 740 1176 1111
+ 1116 583 741 584 1117 1115 742 586 595 1177 743 587 592 744 588 745 746 589 1118 747
+ 1178 748 1179 590 750 591 753 1120 751 749 752 594 759 754 755 756 605 758 597 757
+ 598 610 760 1079 761 602 599 762 600 764 604 763 603 766 765 1016 1181 1137 403 1014
+ 1122 1128 768 1133 611 601 1124 1130 1134 1125 606 1123 607 769 1136 1127 1135 608 770 1139
+ 1185 772 1190 1131 1132 1126 609 771 773 1129 651 1183 774 775 1182 886 612 1184 1138 1186
+ 776 835 613 1187 1188 887 614 777 778 1141 781 615 779 1191 1189 616 617 780 618 782
+ 619 620 784 783 1140 1192 788 786 785 1194 1193 787 621 622 789 1195 623 624 790 791
+ 792 626 793 625 627 794 628 629 795 630 631 632 633 634 636 796 798 797 637 635
+ 799 800 802 801 639 640 803 641 804 1180 643 638 644 642 1142 1143 806 1196 1199 808
+ 646 1144 809 1197 1198 645 1149 1146 1201 648 1200 810 1145 807 805 649 811 1150 812 655
+ 1148 650 813 652 654 885 653 1151 647 658 814 656 657 815 1152 818 816 660 659 661
+ 1153 817 1052 1154 1157 1159 1155 1156 662 664 819 665 666 668 673 1163 667 672 1160 669
+ 670 820 821 1161 671 1162 1168 823 1164 824 680 674 1165 829 822 1158 675 663 825 827
+ 826 676 1169 679 678 828 683 1166 682 1170 681 830 699 684 677 832 831 686 685 12
+ 693 833 1171 1202 687 688 689 834 708 691 692 690 837 836 1172 694 838 695 839 840
+ 841 696 698 697 852 1167 700 1173 843 701 842 1203 702 1174 1 846 844 860 845 868
+ 704 703 511 871 849 1175 707 705 848 847 706 850 709 851 710 853 711 855 854 712
+ 716 713 714 858 725 715 856 857 8 717 718 719 859 720 722 721 724 723 7 67
+ 1222
+ ICV_24 $T=0 0 0 0 $X=139500 $Y=391180
X15 GND VCC 40 38 41 729 734 732 730 731 733 738 737 739 736 1176 740 735 741 742
+ 747 743 1178 744 745 1177 748 749 751 750 1179 752 754 753 755 746 756 757 759 1180
+ 758 760 761 766 763 764 762 765 1181 804 767 803 768 769 1196 1193 771 772 770 1183
+ 1182 773 886 774 1186 1184 775 778 1185 1188 776 777 1189 1190 792 1187 779 1191 780 781
+ 783 784 785 1192 786 1194 787 887 1195 788 789 791 790 782 793 794 1197 795 796 797
+ 798 799 48 800 801 802 809 1199 1201 805 806 810 1198 1200 807 808 813 811 812 816
+ 814 815 817 818 819 824 820 823 49 826 1202 825 828 829 830 832 831 833 836 834
+ 835 867 837 838 839 840 841 1203 852 854 842 843 845 846 847 848 849 850 32 857
+ 851 853 855 858 856 859 67 68 69 1222
+ ICV_25 $T=0 0 0 0 $X=139500 $Y=139500
X16 40 41 48 49 o_data[0] 821 32 o_data[1] 822 o_data[2] 827 o_data[8] 867 868 857 o_data[9] 860 68 i_data[6] 726
+ i_data[7] 727 1222
+ ICV_26 $T=0 0 0 0 $X=139500 $Y=-56920
X18 32 33 o_data[14] 82 879 1222 ICV_28 $T=0 0 0 0 $X=-56920 $Y=1077400
X19 i_data[5] 82 880 1222 ICV_29 $T=0 0 0 0 $X=-56920 $Y=900200
X20 36 i_data[4] 550 1222 ICV_30 $T=0 0 0 0 $X=-56920 $Y=719600
X22 37 36 i_data[3] 1222 ICV_32 $T=0 0 0 0 $X=-56920 $Y=391200
X23 38 39 i_data[1] 728 i_data[2] 1222 ICV_33 $T=0 0 0 0 $X=-56920 $Y=139500
.ENDS
***************************************
